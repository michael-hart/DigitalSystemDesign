LIBRARY IEEE;

USE IEEE.std_logic_1164.ALL;

PACKAGE fp_mult_data_pak IS

	-- Define data types array
	TYPE data_t_rec IS
		RECORD
      		dataa, datab, result : std_logic_vector(31 DOWNTO 0);
		END RECORD;
	TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;
	
	-- Define actual data
	CONSTANT data : data_t := (
		(X"00000000", X"00000000", X"00000000"),
		(X"3dcccccd", X"00000000", X"3d6ef844"),
		(X"3e4ccccd", X"00000000", X"3e0891de"),
		(X"3e99999a", X"00000000", X"3e667b66"),
		(X"3ecccccd", X"00000000", X"3eaabd55"),
		(X"3f000000", X"00000000", X"3eeac7d5"),
		(X"3f19999a", X"00000000", X"3f19ae99"),
		(X"3f333333", X"00000000", X"3f423eb7"),
		(X"3f4ccccd", X"00000000", X"3f6f1444"),
		(X"3f666666", X"00000000", X"3f9017a0"),
		(X"3f800000", X"00000000", X"3faac7d5"),
		(X"3f8ccccd", X"00000000", X"3fc79ac1"),
		(X"3f99999a", X"00000000", X"3fe69066"),
		(X"3fa66666", X"00000000", X"4003d461"),
		(X"3fb33333", X"00000000", X"401571ea"),
		(X"3fc00000", X"00000000", X"402820cf"),
		(X"3fcccccd", X"00000000", X"403be110"),
		(X"3fd9999a", X"00000000", X"4050b2ad"),
		(X"3fe66666", X"00000000", X"406695a5"),
		(X"3ff33333", X"00000000", X"407d89fa"),
		(X"40000000", X"00000000", X"408ac7d5"),
		(X"40066666", X"00000000", X"4097535b"),
		(X"400ccccd", X"00000000", X"40a4678e"),
		(X"40133333", X"00000000", X"40b20470"),
		(X"4019999a", X"00000000", X"40c029ff"),
		(X"40200000", X"00000000", X"40ced83c"),
		(X"40266666", X"00000000", X"40de0f28"),
		(X"402ccccd", X"00000000", X"40edcec1"),
		(X"40333333", X"00000000", X"40fe1707"),
		(X"4039999a", X"00000000", X"410773fe"),
		(X"40400000", X"00000000", X"411020cf"),
		(X"40466666", X"00000000", X"411911f8"),
		(X"404ccccd", X"00000000", X"41224777"),
		(X"40533333", X"00000000", X"412bc14d"),
		(X"4059999a", X"00000000", X"41357f7a"),
		(X"40600000", X"00000000", X"413f81fe"),
		(X"40666666", X"00000000", X"4149c8d9"),
		(X"406ccccd", X"00000000", X"4154540a"),
		(X"40733333", X"00000000", X"415f2393"),
		(X"4079999a", X"00000000", X"416a3773"),
		(X"40800000", X"00000000", X"41851647"),
		(X"40833333", X"00000000", X"418b6a20"),
		(X"40866666", X"00000000", X"4191e371"),
		(X"4089999a", X"00000000", X"41988239"),
		(X"408ccccd", X"00000000", X"419f467a"),
		(X"40900000", X"00000000", X"41a63032"),
		(X"40933333", X"00000000", X"41ad3f62"),
		(X"40966666", X"00000000", X"41b47409"),
		(X"4099999a", X"00000000", X"41bbce29"),
		(X"409ccccd", X"00000000", X"41c34dc0"),
		(X"40a00000", X"00000000", X"41caf2cf"),
		(X"40a33333", X"00000000", X"41d2bd56"),
		(X"40a66666", X"00000000", X"41daad54"),
		(X"40a9999a", X"00000000", X"41e2c2cb"),
		(X"40accccd", X"00000000", X"41eafdb9"),
		(X"40b00000", X"00000000", X"41f35e1e"),
		(X"40b33333", X"00000000", X"41fbe3fc"),
		(X"40b66666", X"00000000", X"420247a9"),
		(X"40b9999a", X"00000000", X"4206b00f"),
		(X"40bccccd", X"00000000", X"420b2b32"),
		(X"40c00000", X"00000000", X"420fb910"),
		(X"40c33333", X"00000000", X"421459aa"),
		(X"40c66666", X"00000000", X"42190d00"),
		(X"40c9999a", X"00000000", X"421dd312"),
		(X"40cccccd", X"00000000", X"4222abe0"),
		(X"40d00000", X"00000000", X"4227976a"),
		(X"40d33333", X"00000000", X"422c95af"),
		(X"40d66666", X"00000000", X"4231a6b1"),
		(X"40d9999a", X"00000000", X"4236ca6e"),
		(X"40dccccd", X"00000000", X"423c00e8"),
		(X"40e00000", X"00000000", X"42414a1d"),
		(X"40e33333", X"00000000", X"4246a60e"),
		(X"40e66666", X"00000000", X"424c14bb"),
		(X"40e9999a", X"00000000", X"42519624"),
		(X"40eccccd", X"00000000", X"42572a48"),
		(X"40f00000", X"00000000", X"425cd129"),
		(X"40f33333", X"00000000", X"42628ac5"),
		(X"40f66666", X"00000000", X"4268571e"),
		(X"40f9999a", X"00000000", X"426e3632"),
		(X"40fccccd", X"00000000", X"42742802"),
		(X"41000000", X"00000000", X"415df418"),
		(X"4101999a", X"00000000", X"4162ba1d"),
		(X"41033333", X"00000000", X"41678cc5"),
		(X"4104cccd", X"00000000", X"416c6c10"),
		(X"41066666", X"00000000", X"417157fe"),
		(X"41080000", X"00000000", X"4176508f"),
		(X"4109999a", X"00000000", X"417b55c2"),
		(X"410b3333", X"00000000", X"418033cc"),
		(X"410ccccd", X"00000000", X"4182c309"),
		(X"410e6666", X"00000000", X"41855897"),
		(X"41100000", X"00000000", X"4187f477"),
		(X"4111999a", X"00000000", X"418a96a8"),
		(X"41133333", X"00000000", X"418d3f2a"),
		(X"4114cccd", X"00000000", X"418fedfe"),
		(X"41166666", X"00000000", X"4192a324"),
		(X"41180000", X"00000000", X"41955e9b"),
		(X"4119999a", X"00000000", X"41982063"),
		(X"411b3333", X"00000000", X"419ae87d"),
		(X"411ccccd", X"00000000", X"419db6e8"),
		(X"411e6666", X"00000000", X"41a08ba4"),
		(X"41200000", X"00000000", X"41a366b2"),
		(X"4121999a", X"00000000", X"41a64812"),
		(X"41233333", X"00000000", X"41a92fc3"),
		(X"4124cccd", X"00000000", X"41ac1dc5"),
		(X"41266666", X"00000000", X"41af1219"),
		(X"41280000", X"00000000", X"41b20cbe"),
		(X"4129999a", X"00000000", X"41b50db5"),
		(X"412b3333", X"00000000", X"41b814fd"),
		(X"412ccccd", X"00000000", X"41bb2297"),
		(X"412e6666", X"00000000", X"41be3682"),
		(X"41300000", X"00000000", X"41c150be"),
		(X"4131999a", X"00000000", X"41c4714c"),
		(X"41333333", X"00000000", X"41c7982c"),
		(X"4134cccd", X"00000000", X"41cac55c"),
		(X"41366666", X"00000000", X"41cdf8df"),
		(X"41380000", X"00000000", X"41d132b2"),
		(X"4139999a", X"00000000", X"41d472d8"),
		(X"413b3333", X"00000000", X"41d7b94e"),
		(X"413ccccd", X"00000000", X"41db0616"),
		(X"413e6666", X"00000000", X"41de5930"),
		(X"41400000", X"00000000", X"c2cb70c9"),
		(X"4141999a", X"00000000", X"c2cef23b"),
		(X"41433333", X"00000000", X"c2d27b55"),
		(X"4144cccd", X"00000000", X"c2d60c18"),
		(X"41466666", X"00000000", X"c2d9a485"),
		(X"41480000", X"00000000", X"c2dd449a"),
		(X"4149999a", X"00000000", X"c2e0ec59"),
		(X"414b3333", X"00000000", X"c2e49bc0"),
		(X"414ccccd", X"00000000", X"c2e852d0"),
		(X"414e6666", X"00000000", X"c2ec118a"),
		(X"41500000", X"00000000", X"c2efd7ec"),
		(X"4151999a", X"00000000", X"c2f3a5f7"),
		(X"41533333", X"00000000", X"c2f77bac"),
		(X"4154cccd", X"00000000", X"c2fb5909"),
		(X"41566666", X"00000000", X"c2ff3e0f"),
		(X"41580000", X"00000000", X"c301955f"),
		(X"4159999a", X"00000000", X"c3038f8b"),
		(X"415b3333", X"00000000", X"c3058d8c"),
		(X"415ccccd", X"00000000", X"c3078f61"),
		(X"415e6666", X"00000000", X"c309950b"),
		(X"41600000", X"00000000", X"c30b9e89"),
		(X"4161999a", X"00000000", X"c30dabdb"),
		(X"41633333", X"00000000", X"c30fbd03"),
		(X"4164cccd", X"00000000", X"c311d1fe"),
		(X"41666666", X"00000000", X"c313eace"),
		(X"41680000", X"00000000", X"c3160773"),
		(X"4169999a", X"00000000", X"c31827ec"),
		(X"416b3333", X"00000000", X"c31a4c39"),
		(X"416ccccd", X"00000000", X"c31c745c"),
		(X"416e6666", X"00000000", X"c31ea052"),
		(X"41700000", X"00000000", X"c320d01d"),
		(X"4171999a", X"00000000", X"c32303bd"),
		(X"41733333", X"00000000", X"c3253b31"),
		(X"4174cccd", X"00000000", X"c3277679"),
		(X"41766666", X"00000000", X"c329b596"),
		(X"41780000", X"00000000", X"c32bf888"),
		(X"4179999a", X"00000000", X"c32e3f4e"),
		(X"417b3333", X"00000000", X"c33089e8"),
		(X"417ccccd", X"00000000", X"c332d857"),
		(X"417e6666", X"00000000", X"c3352a9b"),
		(X"41800000", X"00000000", X"c36e6d57"),
		(X"4180cccd", X"00000000", X"c3717792"),
		(X"4181999a", X"00000000", X"c37486bb"),
		(X"41826666", X"00000000", X"c3779ad1"),
		(X"41833333", X"00000000", X"c37ab3d5"),
		(X"41840000", X"00000000", X"c37dd1c7"),
		(X"4184cccd", X"00000000", X"c3807a53"),
		(X"4185999a", X"00000000", X"c3820e3a"),
		(X"41866666", X"00000000", X"c383a498"),
		(X"41873333", X"00000000", X"c3853d6c"),
		(X"41880000", X"00000000", X"c386d8b7"),
		(X"4188cccd", X"00000000", X"c3887679"),
		(X"4189999a", X"00000000", X"c38a16b2"),
		(X"418a6666", X"00000000", X"c38bb962"),
		(X"418b3333", X"00000000", X"c38d5e89"),
		(X"418c0000", X"00000000", X"c38f0626"),
		(X"418ccccd", X"00000000", X"c390b03b"),
		(X"418d999a", X"00000000", X"c3925cc6"),
		(X"418e6666", X"00000000", X"c3940bc8"),
		(X"418f3333", X"00000000", X"c395bd41"),
		(X"41900000", X"00000000", X"c3977131"),
		(X"4190cccd", X"00000000", X"c3992797"),
		(X"4191999a", X"00000000", X"c39ae075"),
		(X"41926666", X"00000000", X"c39c9bc9"),
		(X"41933333", X"00000000", X"c39e5994"),
		(X"41940000", X"00000000", X"c3a019d6"),
		(X"4194cccd", X"00000000", X"c3a1dc8f"),
		(X"4195999a", X"00000000", X"c3a3a1bf"),
		(X"41966666", X"00000000", X"c3a56966"),
		(X"41973333", X"00000000", X"c3a73383"),
		(X"41980000", X"00000000", X"c3a90018"),
		(X"4198cccd", X"00000000", X"c3aacf23"),
		(X"4199999a", X"00000000", X"c3aca0a5"),
		(X"419a6666", X"00000000", X"c3ae749e"),
		(X"419b3333", X"00000000", X"c3b04b0d"),
		(X"419c0000", X"00000000", X"c3b223f4"),
		(X"419ccccd", X"00000000", X"c3b3ff51"),
		(X"419d999a", X"00000000", X"c3b5dd26"),
		(X"419e6666", X"00000000", X"c3b7bd71"),
		(X"419f3333", X"00000000", X"c3b9a033"),
		(X"41a00000", X"00000000", X"c2d5b607"),
		(X"41a0cccd", X"00000000", X"c2d7f439"),
		(X"41a1999a", X"00000000", X"c2da3569"),
		(X"41a26666", X"00000000", X"c2dc7997"),
		(X"41a33333", X"00000000", X"c2dec0c3"),
		(X"41a40000", X"00000000", X"c2e10aec"),
		(X"41a4cccd", X"00000000", X"c2e35814"),
		(X"41a5999a", X"00000000", X"c2e5a839"),
		(X"41a66666", X"00000000", X"c2e7fb5c"),
		(X"41a73333", X"00000000", X"c2ea517d"),
		(X"41a80000", X"00000000", X"c2ecaa9b"),
		(X"41a8cccd", X"00000000", X"c2ef06b8"),
		(X"41a9999a", X"00000000", X"c2f165d2"),
		(X"41aa6666", X"00000000", X"c2f3c7ea"),
		(X"41ab3333", X"00000000", X"c2f62d00"),
		(X"41ac0000", X"00000000", X"c2f89513"),
		(X"41accccd", X"00000000", X"c2fb0025"),
		(X"41ad999a", X"00000000", X"c2fd6e34"),
		(X"41ae6666", X"00000000", X"c2ffdf42"),
		(X"41af3333", X"00000000", X"c30129a6"),
		(X"41b00000", X"00000000", X"c302652b"),
		(X"41b0cccd", X"00000000", X"c303a22e"),
		(X"41b1999a", X"00000000", X"c304e0b0"),
		(X"41b26666", X"00000000", X"c30620b1"),
		(X"41b33333", X"00000000", X"c3076232"),
		(X"41b40000", X"00000000", X"c308a531"),
		(X"41b4cccd", X"00000000", X"c309e9ae"),
		(X"41b5999a", X"00000000", X"c30b2fab"),
		(X"41b66666", X"00000000", X"c30c7727"),
		(X"41b73333", X"00000000", X"c30dc022"),
		(X"41b80000", X"00000000", X"c30f0a9b"),
		(X"41b8cccd", X"00000000", X"c3105694"),
		(X"41b9999a", X"00000000", X"c311a40b"),
		(X"41ba6666", X"00000000", X"c312f301"),
		(X"41bb3333", X"00000000", X"c3144376"),
		(X"41bc0000", X"00000000", X"c315956b"),
		(X"41bccccd", X"00000000", X"c316e8de"),
		(X"41bd999a", X"00000000", X"c3183dd0"),
		(X"41be6666", X"00000000", X"c3199440"),
		(X"41bf3333", X"00000000", X"c31aec30"),
		(X"41c00000", X"00000000", X"43c05011"),
		(X"41c0cccd", X"00000000", X"43c1e4c3"),
		(X"41c1999a", X"00000000", X"43c37b1d"),
		(X"41c26666", X"00000000", X"43c5131f"),
		(X"41c33333", X"00000000", X"43c6acc9"),
		(X"41c40000", X"00000000", X"43c8481b"),
		(X"41c4cccd", X"00000000", X"43c9e515"),
		(X"41c5999a", X"00000000", X"43cb83b7"),
		(X"41c66666", X"00000000", X"43cd2400"),
		(X"41c73333", X"00000000", X"43cec5f2"),
		(X"41c80000", X"00000000", X"43d0698c"),
		(X"41c8cccd", X"00000000", X"43d20ecd"),
		(X"41c9999a", X"00000000", X"43d3b5b7"),
		(X"41ca6666", X"00000000", X"43d55e49"),
		(X"41cb3333", X"00000000", X"43d70882"),
		(X"41cc0000", X"00000000", X"43d8b464"),
		(X"41cccccd", X"00000000", X"43da61ed"),
		(X"41cd999a", X"00000000", X"43dc111e"),
		(X"41ce6666", X"00000000", X"43ddc1f8"),
		(X"41cf3333", X"00000000", X"43df7479"),
		(X"41d00000", X"00000000", X"43e128a3"),
		(X"41d0cccd", X"00000000", X"43e2de74"),
		(X"41d1999a", X"00000000", X"43e495ed"),
		(X"41d26666", X"00000000", X"43e64f0e"),
		(X"41d33333", X"00000000", X"43e809d8"),
		(X"41d40000", X"00000000", X"43e9c649"),
		(X"41d4cccd", X"00000000", X"43eb8462"),
		(X"41d5999a", X"00000000", X"43ed4423"),
		(X"41d66666", X"00000000", X"43ef058c"),
		(X"41d73333", X"00000000", X"43f0c89d"),
		(X"41d80000", X"00000000", X"43f28d56"),
		(X"41d8cccd", X"00000000", X"43f453b7"),
		(X"41d9999a", X"00000000", X"43f61bc0"),
		(X"41da6666", X"00000000", X"43f7e571"),
		(X"41db3333", X"00000000", X"43f9b0ca"),
		(X"41dc0000", X"00000000", X"43fb7dca"),
		(X"41dccccd", X"00000000", X"43fd4c73"),
		(X"41dd999a", X"00000000", X"43ff1cc4"),
		(X"41de6666", X"00000000", X"4400775e"),
		(X"41df3333", X"00000000", X"4401612f"),
		(X"41e00000", X"00000000", X"4445c698"),
		(X"41e0cccd", X"00000000", X"44472dac"),
		(X"41e1999a", X"00000000", X"44489606"),
		(X"41e26666", X"00000000", X"4449ffa5"),
		(X"41e33333", X"00000000", X"444b6a88"),
		(X"41e40000", X"00000000", X"444cd6b0"),
		(X"41e4cccd", X"00000000", X"444e441d"),
		(X"41e5999a", X"00000000", X"444fb2ce"),
		(X"41e66666", X"00000000", X"445122c5"),
		(X"41e73333", X"00000000", X"44529400"),
		(X"41e80000", X"00000000", X"44540680"),
		(X"41e8cccd", X"00000000", X"44557a45"),
		(X"41e9999a", X"00000000", X"4456ef4e"),
		(X"41ea6666", X"00000000", X"4458659d"),
		(X"41eb3333", X"00000000", X"4459dd30"),
		(X"41ec0000", X"00000000", X"445b5608"),
		(X"41eccccd", X"00000000", X"445cd025"),
		(X"41ed999a", X"00000000", X"445e4b87"),
		(X"41ee6666", X"00000000", X"445fc82d"),
		(X"41ef3333", X"00000000", X"44614618"),
		(X"41f00000", X"00000000", X"4462c548"),
		(X"41f0cccd", X"00000000", X"446445bd"),
		(X"41f1999a", X"00000000", X"4465c777"),
		(X"41f26666", X"00000000", X"44674a75"),
		(X"41f33333", X"00000000", X"4468ceb8"),
		(X"41f40000", X"00000000", X"446a5440"),
		(X"41f4cccd", X"00000000", X"446bdb0d"),
		(X"41f5999a", X"00000000", X"446d631f"),
		(X"41f66666", X"00000000", X"446eec75"),
		(X"41f73333", X"00000000", X"44707710"),
		(X"41f80000", X"00000000", X"447202f0"),
		(X"41f8cccd", X"00000000", X"44739015"),
		(X"41f9999a", X"00000000", X"44751e7e"),
		(X"41fa6666", X"00000000", X"4476ae2d"),
		(X"41fb3333", X"00000000", X"44783f20"),
		(X"41fc0000", X"00000000", X"4479d158"),
		(X"41fccccd", X"00000000", X"447b64d5"),
		(X"41fd999a", X"00000000", X"447cf996"),
		(X"41fe6666", X"00000000", X"447e8f9d"),
		(X"41ff3333", X"00000000", X"44801374"),
		(X"42000000", X"00000000", X"43e12dfe"),
		(X"42006666", X"00000000", X"43e2906c"),
		(X"4200cccd", X"00000000", X"43e3f3f0"),
		(X"42013333", X"00000000", X"43e5588a"),
		(X"4201999a", X"00000000", X"43e6be3a"),
		(X"42020000", X"00000000", X"43e82500"),
		(X"42026666", X"00000000", X"43e98cdd"),
		(X"4202cccd", X"00000000", X"43eaf5cf"),
		(X"42033333", X"00000000", X"43ec5fd7"),
		(X"4203999a", X"00000000", X"43edcaf5"),
		(X"42040000", X"00000000", X"43ef3729"),
		(X"42046666", X"00000000", X"43f0a473"),
		(X"4204cccd", X"00000000", X"43f212d3"),
		(X"42053333", X"00000000", X"43f38249"),
		(X"4205999a", X"00000000", X"43f4f2d5"),
		(X"42060000", X"00000000", X"43f66477"),
		(X"42066666", X"00000000", X"43f7d72f"),
		(X"4206cccd", X"00000000", X"43f94afd"),
		(X"42073333", X"00000000", X"43fabfe1"),
		(X"4207999a", X"00000000", X"43fc35db"),
		(X"42080000", X"00000000", X"43fdaceb"),
		(X"42086666", X"00000000", X"43ff2511"),
		(X"4208cccd", X"00000000", X"44004f27"),
		(X"42093333", X"00000000", X"44010c50"),
		(X"4209999a", X"00000000", X"4401ca04"),
		(X"420a0000", X"00000000", X"44028843"),
		(X"420a6666", X"00000000", X"4403470d"),
		(X"420acccd", X"00000000", X"44040662"),
		(X"420b3333", X"00000000", X"4404c641"),
		(X"420b999a", X"00000000", X"440586ac"),
		(X"420c0000", X"00000000", X"440647a2"),
		(X"420c6666", X"00000000", X"44070923"),
		(X"420ccccd", X"00000000", X"4407cb2f"),
		(X"420d3333", X"00000000", X"44088dc6"),
		(X"420d999a", X"00000000", X"440950e8"),
		(X"420e0000", X"00000000", X"440a1495"),
		(X"420e6666", X"00000000", X"440ad8cd"),
		(X"420ecccd", X"00000000", X"440b9d90"),
		(X"420f3333", X"00000000", X"440c62de"),
		(X"420f999a", X"00000000", X"440d28b7"),
		(X"42100000", X"00000000", X"c428234d"),
		(X"42106666", X"00000000", X"c42915f9"),
		(X"4210cccd", X"00000000", X"c42a0953"),
		(X"42113333", X"00000000", X"c42afd5c"),
		(X"4211999a", X"00000000", X"c42bf213"),
		(X"42120000", X"00000000", X"c42ce77a"),
		(X"42126666", X"00000000", X"c42ddd8e"),
		(X"4212cccd", X"00000000", X"c42ed451"),
		(X"42133333", X"00000000", X"c42fcbc3"),
		(X"4213999a", X"00000000", X"c430c3e4"),
		(X"42140000", X"00000000", X"c431bcb3"),
		(X"42146666", X"00000000", X"c432b630"),
		(X"4214cccd", X"00000000", X"c433b05d"),
		(X"42153333", X"00000000", X"c434ab37"),
		(X"4215999a", X"00000000", X"c435a6c1"),
		(X"42160000", X"00000000", X"c436a2f9"),
		(X"42166666", X"00000000", X"c4379fdf"),
		(X"4216cccd", X"00000000", X"c4389d75"),
		(X"42173333", X"00000000", X"c4399bb8"),
		(X"4217999a", X"00000000", X"c43a9aab"),
		(X"42180000", X"00000000", X"c43b9a4c"),
		(X"42186666", X"00000000", X"c43c9a9b"),
		(X"4218cccd", X"00000000", X"c43d9b9a"),
		(X"42193333", X"00000000", X"c43e9d47"),
		(X"4219999a", X"00000000", X"c43f9fa2"),
		(X"421a0000", X"00000000", X"c440a2ac"),
		(X"421a6666", X"00000000", X"c441a665"),
		(X"421acccd", X"00000000", X"c442aacc"),
		(X"421b3333", X"00000000", X"c443afe2"),
		(X"421b999a", X"00000000", X"c444b5a6"),
		(X"421c0000", X"00000000", X"c445bc19"),
		(X"421c6666", X"00000000", X"c446c33b"),
		(X"421ccccd", X"00000000", X"c447cb0b"),
		(X"421d3333", X"00000000", X"c448d38a"),
		(X"421d999a", X"00000000", X"c449dcb7"),
		(X"421e0000", X"00000000", X"c44ae693"),
		(X"421e6666", X"00000000", X"c44bf11e"),
		(X"421ecccd", X"00000000", X"c44cfc57"),
		(X"421f3333", X"00000000", X"c44e083f"),
		(X"421f999a", X"00000000", X"c44f14d5"),
		(X"42200000", X"00000000", X"c4c57dff"),
		(X"42206666", X"00000000", X"c4c67cb4"),
		(X"4220cccd", X"00000000", X"c4c77c0e"),
		(X"42213333", X"00000000", X"c4c87c0b"),
		(X"4221999a", X"00000000", X"c4c97cad"),
		(X"42220000", X"00000000", X"c4ca7df2"),
		(X"42226666", X"00000000", X"c4cb7fdb"),
		(X"4222cccd", X"00000000", X"c4cc8267"),
		(X"42233333", X"00000000", X"c4cd8598"),
		(X"4223999a", X"00000000", X"c4ce896c"),
		(X"42240000", X"00000000", X"c4cf8de5"),
		(X"42246666", X"00000000", X"c4d09301"),
		(X"4224cccd", X"00000000", X"c4d198c1"),
		(X"42253333", X"00000000", X"c4d29f24"),
		(X"4225999a", X"00000000", X"c4d3a62c"),
		(X"42260000", X"00000000", X"c4d4add7"),
		(X"42266666", X"00000000", X"c4d5b627"),
		(X"4226cccd", X"00000000", X"c4d6bf1a"),
		(X"42273333", X"00000000", X"c4d7c8b1"),
		(X"4227999a", X"00000000", X"c4d8d2eb"),
		(X"42280000", X"00000000", X"c4d9ddca"),
		(X"42286666", X"00000000", X"c4dae94c"),
		(X"4228cccd", X"00000000", X"c4dbf573"),
		(X"42293333", X"00000000", X"c4dd023d"),
		(X"4229999a", X"00000000", X"c4de0fab"),
		(X"422a0000", X"00000000", X"c4df1dbc"),
		(X"422a6666", X"00000000", X"c4e02c72"),
		(X"422acccd", X"00000000", X"c4e13bcb"),
		(X"422b3333", X"00000000", X"c4e24bc9"),
		(X"422b999a", X"00000000", X"c4e35c6a"),
		(X"422c0000", X"00000000", X"c4e46daf"),
		(X"422c6666", X"00000000", X"c4e57f97"),
		(X"422ccccd", X"00000000", X"c4e69224"),
		(X"422d3333", X"00000000", X"c4e7a554"),
		(X"422d999a", X"00000000", X"c4e8b929"),
		(X"422e0000", X"00000000", X"c4e9cda1"),
		(X"422e6666", X"00000000", X"c4eae2bd"),
		(X"422ecccd", X"00000000", X"c4ebf87c"),
		(X"422f3333", X"00000000", X"c4ed0ee0"),
		(X"422f999a", X"00000000", X"c4ee25e7"),
		(X"42300000", X"00000000", X"c481ccec"),
		(X"42306666", X"00000000", X"c48265bd"),
		(X"4230cccd", X"00000000", X"c482fee8"),
		(X"42313333", X"00000000", X"c483986c"),
		(X"4231999a", X"00000000", X"c484324a"),
		(X"42320000", X"00000000", X"c484cc82"),
		(X"42326666", X"00000000", X"c4856714"),
		(X"4232cccd", X"00000000", X"c48601ff"),
		(X"42333333", X"00000000", X"c4869d44"),
		(X"4233999a", X"00000000", X"c48738e3"),
		(X"42340000", X"00000000", X"c487d4db"),
		(X"42346666", X"00000000", X"c488712d"),
		(X"4234cccd", X"00000000", X"c4890dd9"),
		(X"42353333", X"00000000", X"c489aadf"),
		(X"4235999a", X"00000000", X"c48a483f"),
		(X"42360000", X"00000000", X"c48ae5f8"),
		(X"42366666", X"00000000", X"c48b840b"),
		(X"4236cccd", X"00000000", X"c48c2277"),
		(X"42373333", X"00000000", X"c48cc13e"),
		(X"4237999a", X"00000000", X"c48d605e"),
		(X"42380000", X"00000000", X"c48dffd8"),
		(X"42386666", X"00000000", X"c48e9fac"),
		(X"4238cccd", X"00000000", X"c48f3fd9"),
		(X"42393333", X"00000000", X"c48fe060"),
		(X"4239999a", X"00000000", X"c4908141"),
		(X"423a0000", X"00000000", X"c491227c"),
		(X"423a6666", X"00000000", X"c491c410"),
		(X"423acccd", X"00000000", X"c49265fe"),
		(X"423b3333", X"00000000", X"c4930846"),
		(X"423b999a", X"00000000", X"c493aae7"),
		(X"423c0000", X"00000000", X"c4944de3"),
		(X"423c6666", X"00000000", X"c494f138"),
		(X"423ccccd", X"00000000", X"c49594e7"),
		(X"423d3333", X"00000000", X"c49638ef"),
		(X"423d999a", X"00000000", X"c496dd51"),
		(X"423e0000", X"00000000", X"c497820d"),
		(X"423e6666", X"00000000", X"c4982723"),
		(X"423ecccd", X"00000000", X"c498cc93"),
		(X"423f3333", X"00000000", X"c499725c"),
		(X"423f999a", X"00000000", X"c49a187f"),
		(X"42400000", X"00000000", X"44710e26"),
		(X"42406666", X"00000000", X"44720c56"),
		(X"4240cccd", X"00000000", X"44730b0b"),
		(X"42413333", X"00000000", X"44740a47"),
		(X"4241999a", X"00000000", X"44750a08"),
		(X"42420000", X"00000000", X"44760a4e"),
		(X"42426666", X"00000000", X"44770b1b"),
		(X"4242cccd", X"00000000", X"44780c6d"),
		(X"42433333", X"00000000", X"44790e45"),
		(X"4243999a", X"00000000", X"447a10a2"),
		(X"42440000", X"00000000", X"447b1386"),
		(X"42446666", X"00000000", X"447c16ef"),
		(X"4244cccd", X"00000000", X"447d1add"),
		(X"42453333", X"00000000", X"447e1f52"),
		(X"4245999a", X"00000000", X"447f244c"),
		(X"42460000", X"00000000", X"448014e6"),
		(X"42466666", X"00000000", X"448097e9"),
		(X"4246cccd", X"00000000", X"44811b2e"),
		(X"42473333", X"00000000", X"44819eb7"),
		(X"4247999a", X"00000000", X"44822282"),
		(X"42480000", X"00000000", X"4482a691"),
		(X"42486666", X"00000000", X"44832ae2"),
		(X"4248cccd", X"00000000", X"4483af76"),
		(X"42493333", X"00000000", X"4484344d"),
		(X"4249999a", X"00000000", X"4484b966"),
		(X"424a0000", X"00000000", X"44853ec3"),
		(X"424a6666", X"00000000", X"4485c462"),
		(X"424acccd", X"00000000", X"44864a44"),
		(X"424b3333", X"00000000", X"4486d06a"),
		(X"424b999a", X"00000000", X"448756d2"),
		(X"424c0000", X"00000000", X"4487dd7c"),
		(X"424c6666", X"00000000", X"4488646a"),
		(X"424ccccd", X"00000000", X"4488eb9b"),
		(X"424d3333", X"00000000", X"4489730e"),
		(X"424d999a", X"00000000", X"4489fac4"),
		(X"424e0000", X"00000000", X"448a82be"),
		(X"424e6666", X"00000000", X"448b0afa"),
		(X"424ecccd", X"00000000", X"448b9379"),
		(X"424f3333", X"00000000", X"448c1c3a"),
		(X"424f999a", X"00000000", X"448ca53f"),
		(X"42500000", X"00000000", X"4528b751"),
		(X"42506666", X"00000000", X"45295ccc"),
		(X"4250cccd", X"00000000", X"452a0297"),
		(X"42513333", X"00000000", X"452aa8b4"),
		(X"4251999a", X"00000000", X"452b4f21"),
		(X"42520000", X"00000000", X"452bf5e0"),
		(X"42526666", X"00000000", X"452c9cef"),
		(X"4252cccd", X"00000000", X"452d4450"),
		(X"42533333", X"00000000", X"452dec01"),
		(X"4253999a", X"00000000", X"452e9404"),
		(X"42540000", X"00000000", X"452f3c57"),
		(X"42546666", X"00000000", X"452fe4fc"),
		(X"4254cccd", X"00000000", X"45308df1"),
		(X"42553333", X"00000000", X"45313738"),
		(X"4255999a", X"00000000", X"4531e0cf"),
		(X"42560000", X"00000000", X"45328ab7"),
		(X"42566666", X"00000000", X"453334f1"),
		(X"4256cccd", X"00000000", X"4533df7b"),
		(X"42573333", X"00000000", X"45348a57"),
		(X"4257999a", X"00000000", X"45353583"),
		(X"42580000", X"00000000", X"4535e101"),
		(X"42586666", X"00000000", X"45368ccf"),
		(X"4258cccd", X"00000000", X"453738ef"),
		(X"42593333", X"00000000", X"4537e55f"),
		(X"4259999a", X"00000000", X"45389220"),
		(X"425a0000", X"00000000", X"45393f33"),
		(X"425a6666", X"00000000", X"4539ec96"),
		(X"425acccd", X"00000000", X"453a9a4b"),
		(X"425b3333", X"00000000", X"453b4850"),
		(X"425b999a", X"00000000", X"453bf6a6"),
		(X"425c0000", X"00000000", X"453ca54e"),
		(X"425c6666", X"00000000", X"453d5446"),
		(X"425ccccd", X"00000000", X"453e038f"),
		(X"425d3333", X"00000000", X"453eb32a"),
		(X"425d999a", X"00000000", X"453f6315"),
		(X"425e0000", X"00000000", X"45401352"),
		(X"425e6666", X"00000000", X"4540c3df"),
		(X"425ecccd", X"00000000", X"454174bd"),
		(X"425f3333", X"00000000", X"454225ed"),
		(X"425f999a", X"00000000", X"4542d76d"),
		(X"42600000", X"00000000", X"45032c0d"),
		(X"42606666", X"00000000", X"4503a349"),
		(X"4260cccd", X"00000000", X"45041abb"),
		(X"42613333", X"00000000", X"45049263"),
		(X"4261999a", X"00000000", X"45050a42"),
		(X"42620000", X"00000000", X"45058256"),
		(X"42626666", X"00000000", X"4505faa1"),
		(X"4262cccd", X"00000000", X"45067321"),
		(X"42633333", X"00000000", X"4506ebd8"),
		(X"4263999a", X"00000000", X"450764c5"),
		(X"42640000", X"00000000", X"4507dde7"),
		(X"42646666", X"00000000", X"45085740"),
		(X"4264cccd", X"00000000", X"4508d0cf"),
		(X"42653333", X"00000000", X"45094a94"),
		(X"4265999a", X"00000000", X"4509c490"),
		(X"42660000", X"00000000", X"450a3ec1"),
		(X"42666666", X"00000000", X"450ab928"),
		(X"4266cccd", X"00000000", X"450b33c6"),
		(X"42673333", X"00000000", X"450bae99"),
		(X"4267999a", X"00000000", X"450c29a3"),
		(X"42680000", X"00000000", X"450ca4e3"),
		(X"42686666", X"00000000", X"450d2059"),
		(X"4268cccd", X"00000000", X"450d9c05"),
		(X"42693333", X"00000000", X"450e17e7"),
		(X"4269999a", X"00000000", X"450e93ff"),
		(X"426a0000", X"00000000", X"450f104d"),
		(X"426a6666", X"00000000", X"450f8cd2"),
		(X"426acccd", X"00000000", X"4510098c"),
		(X"426b3333", X"00000000", X"4510867d"),
		(X"426b999a", X"00000000", X"451103a3"),
		(X"426c0000", X"00000000", X"45118100"),
		(X"426c6666", X"00000000", X"4511fe93"),
		(X"426ccccd", X"00000000", X"45127c5c"),
		(X"426d3333", X"00000000", X"4512fa5b"),
		(X"426d999a", X"00000000", X"45137890"),
		(X"426e0000", X"00000000", X"4513f6fb"),
		(X"426e6666", X"00000000", X"4514759c"),
		(X"426ecccd", X"00000000", X"4514f473"),
		(X"426f3333", X"00000000", X"45157381"),
		(X"426f999a", X"00000000", X"4515f2c4"),
		(X"42700000", X"00000000", X"c47025a2"),
		(X"42706666", X"00000000", X"c470f5ef"),
		(X"4270cccd", X"00000000", X"c471c697"),
		(X"42713333", X"00000000", X"c4729798"),
		(X"4271999a", X"00000000", X"c47368f4"),
		(X"42720000", X"00000000", X"c4743aaa"),
		(X"42726666", X"00000000", X"c4750cba"),
		(X"4272cccd", X"00000000", X"c475df24"),
		(X"42733333", X"00000000", X"c476b1e8"),
		(X"4273999a", X"00000000", X"c4778507"),
		(X"42740000", X"00000000", X"c478587f"),
		(X"42746666", X"00000000", X"c4792c52"),
		(X"4274cccd", X"00000000", X"c47a007f"),
		(X"42753333", X"00000000", X"c47ad507"),
		(X"4275999a", X"00000000", X"c47ba9e8"),
		(X"42760000", X"00000000", X"c47c7f23"),
		(X"42766666", X"00000000", X"c47d54b9"),
		(X"4276cccd", X"00000000", X"c47e2aa9"),
		(X"42773333", X"00000000", X"c47f00f3"),
		(X"4277999a", X"00000000", X"c47fd797"),
		(X"42780000", X"00000000", X"c480574b"),
		(X"42786666", X"00000000", X"c480c2f7"),
		(X"4278cccd", X"00000000", X"c4812ed0"),
		(X"42793333", X"00000000", X"c4819ad7"),
		(X"4279999a", X"00000000", X"c482070a"),
		(X"427a0000", X"00000000", X"c482736b"),
		(X"427a6666", X"00000000", X"c482dff8"),
		(X"427acccd", X"00000000", X"c4834cb3"),
		(X"427b3333", X"00000000", X"c483b99b"),
		(X"427b999a", X"00000000", X"c48426b0"),
		(X"427c0000", X"00000000", X"c48493f2"),
		(X"427c6666", X"00000000", X"c4850161"),
		(X"427ccccd", X"00000000", X"c4856efd"),
		(X"427d3333", X"00000000", X"c485dcc6"),
		(X"427d999a", X"00000000", X"c4864abd"),
		(X"427e0000", X"00000000", X"c486b8e0"),
		(X"427e6666", X"00000000", X"c4872731"),
		(X"427ecccd", X"00000000", X"c48795ae"),
		(X"427f3333", X"00000000", X"c4880459"),
		(X"427f999a", X"00000000", X"c4887331"),
		(X"42800000", X"00000000", X"c573292c"),
		(X"42803333", X"00000000", X"c573eca7"),
		(X"42806666", X"00000000", X"c574b071"),
		(X"4280999a", X"00000000", X"c5757489"),
		(X"4280cccd", X"00000000", X"c57638f0"),
		(X"42810000", X"00000000", X"c576fda5"),
		(X"42813333", X"00000000", X"c577c2a9"),
		(X"42816666", X"00000000", X"c57887fb"),
		(X"4281999a", X"00000000", X"c5794d9c"),
		(X"4281cccd", X"00000000", X"c57a138a"),
		(X"42820000", X"00000000", X"c57ad9c8"),
		(X"42823333", X"00000000", X"c57ba054"),
		(X"42826666", X"00000000", X"c57c672e"),
		(X"4282999a", X"00000000", X"c57d2e57"),
		(X"4282cccd", X"00000000", X"c57df5ce"),
		(X"42830000", X"00000000", X"c57ebd94"),
		(X"42833333", X"00000000", X"c57f85a8"),
		(X"42836666", X"00000000", X"c5802705"),
		(X"4283999a", X"00000000", X"c5808b5e"),
		(X"4283cccd", X"00000000", X"c580efde"),
		(X"42840000", X"00000000", X"c5815484"),
		(X"42843333", X"00000000", X"c581b953"),
		(X"42846666", X"00000000", X"c5821e48"),
		(X"4284999a", X"00000000", X"c5828365"),
		(X"4284cccd", X"00000000", X"c582e8a9"),
		(X"42850000", X"00000000", X"c5834e14"),
		(X"42853333", X"00000000", X"c583b3a6"),
		(X"42856666", X"00000000", X"c5841960"),
		(X"4285999a", X"00000000", X"c5847f40"),
		(X"4285cccd", X"00000000", X"c584e548"),
		(X"42860000", X"00000000", X"c5854b78"),
		(X"42863333", X"00000000", X"c585b1ce"),
		(X"42866666", X"00000000", X"c586184c"),
		(X"4286999a", X"00000000", X"c5867ef1"),
		(X"4286cccd", X"00000000", X"c586e5bd"),
		(X"42870000", X"00000000", X"c5874cb0"),
		(X"42873333", X"00000000", X"c587b3cb"),
		(X"42876666", X"00000000", X"c5881b0d"),
		(X"4287999a", X"00000000", X"c5888276"),
		(X"4287cccd", X"00000000", X"c588ea06"),
		(X"42880000", X"00000000", X"c5596cc0"),
		(X"42883333", X"00000000", X"c55a1161"),
		(X"42886666", X"00000000", X"c55ab641"),
		(X"4288999a", X"00000000", X"c55b5b5e"),
		(X"4288cccd", X"00000000", X"c55c00ba"),
		(X"42890000", X"00000000", X"c55ca654"),
		(X"42893333", X"00000000", X"c55d4c2d"),
		(X"42896666", X"00000000", X"c55df243"),
		(X"4289999a", X"00000000", X"c55e9898"),
		(X"4289cccd", X"00000000", X"c55f3f2b"),
		(X"428a0000", X"00000000", X"c55fe5fd"),
		(X"428a3333", X"00000000", X"c5608d0c"),
		(X"428a6666", X"00000000", X"c561345a"),
		(X"428a999a", X"00000000", X"c561dbe6"),
		(X"428acccd", X"00000000", X"c56283b0"),
		(X"428b0000", X"00000000", X"c5632bb8"),
		(X"428b3333", X"00000000", X"c563d3ff"),
		(X"428b6666", X"00000000", X"c5647c84"),
		(X"428b999a", X"00000000", X"c5652547"),
		(X"428bcccd", X"00000000", X"c565ce49"),
		(X"428c0000", X"00000000", X"c5667788"),
		(X"428c3333", X"00000000", X"c5672106"),
		(X"428c6666", X"00000000", X"c567cac2"),
		(X"428c999a", X"00000000", X"c56874bd"),
		(X"428ccccd", X"00000000", X"c5691ef5"),
		(X"428d0000", X"00000000", X"c569c96c"),
		(X"428d3333", X"00000000", X"c56a7421"),
		(X"428d6666", X"00000000", X"c56b1f14"),
		(X"428d999a", X"00000000", X"c56bca46"),
		(X"428dcccd", X"00000000", X"c56c75b5"),
		(X"428e0000", X"00000000", X"c56d2163"),
		(X"428e3333", X"00000000", X"c56dcd50"),
		(X"428e6666", X"00000000", X"c56e797a"),
		(X"428e999a", X"00000000", X"c56f25e3"),
		(X"428ecccd", X"00000000", X"c56fd28a"),
		(X"428f0000", X"00000000", X"c5707f6f"),
		(X"428f3333", X"00000000", X"c5712c92"),
		(X"428f6666", X"00000000", X"c571d9f4"),
		(X"428f999a", X"00000000", X"c5728794"),
		(X"428fcccd", X"00000000", X"c5733572"),
		(X"42900000", X"00000000", X"443a3621"),
		(X"42903333", X"00000000", X"443ab76f"),
		(X"42906666", X"00000000", X"443b38e9"),
		(X"4290999a", X"00000000", X"443bba91"),
		(X"4290cccd", X"00000000", X"443c3c65"),
		(X"42910000", X"00000000", X"443cbe66"),
		(X"42913333", X"00000000", X"443d4094"),
		(X"42916666", X"00000000", X"443dc2ef"),
		(X"4291999a", X"00000000", X"443e4577"),
		(X"4291cccd", X"00000000", X"443ec82b"),
		(X"42920000", X"00000000", X"443f4b0c"),
		(X"42923333", X"00000000", X"443fce1a"),
		(X"42926666", X"00000000", X"44405155"),
		(X"4292999a", X"00000000", X"4440d4bd"),
		(X"4292cccd", X"00000000", X"44415851"),
		(X"42930000", X"00000000", X"4441dc13"),
		(X"42933333", X"00000000", X"44426001"),
		(X"42936666", X"00000000", X"4442e41c"),
		(X"4293999a", X"00000000", X"44436863"),
		(X"4293cccd", X"00000000", X"4443ecd8"),
		(X"42940000", X"00000000", X"44447179"),
		(X"42943333", X"00000000", X"4444f647"),
		(X"42946666", X"00000000", X"44457b42"),
		(X"4294999a", X"00000000", X"4446006a"),
		(X"4294cccd", X"00000000", X"444685be"),
		(X"42950000", X"00000000", X"44470b3f"),
		(X"42953333", X"00000000", X"444790ee"),
		(X"42956666", X"00000000", X"444816c8"),
		(X"4295999a", X"00000000", X"44489cd0"),
		(X"4295cccd", X"00000000", X"44492305"),
		(X"42960000", X"00000000", X"4449a966"),
		(X"42963333", X"00000000", X"444a2ff4"),
		(X"42966666", X"00000000", X"444ab6af"),
		(X"4296999a", X"00000000", X"444b3d97"),
		(X"4296cccd", X"00000000", X"444bc4ab"),
		(X"42970000", X"00000000", X"444c4bed"),
		(X"42973333", X"00000000", X"444cd35b"),
		(X"42976666", X"00000000", X"444d5af6"),
		(X"4297999a", X"00000000", X"444de2be"),
		(X"4297cccd", X"00000000", X"444e6ab2"),
		(X"42980000", X"00000000", X"45a4fb4d"),
		(X"42983333", X"00000000", X"45a56a1e"),
		(X"42986666", X"00000000", X"45a5d915"),
		(X"4298999a", X"00000000", X"45a64831"),
		(X"4298cccd", X"00000000", X"45a6b772"),
		(X"42990000", X"00000000", X"45a726d8"),
		(X"42993333", X"00000000", X"45a79663"),
		(X"42996666", X"00000000", X"45a80614"),
		(X"4299999a", X"00000000", X"45a875e9"),
		(X"4299cccd", X"00000000", X"45a8e5e4"),
		(X"429a0000", X"00000000", X"45a95604"),
		(X"429a3333", X"00000000", X"45a9c649"),
		(X"429a6666", X"00000000", X"45aa36b3"),
		(X"429a999a", X"00000000", X"45aaa743"),
		(X"429acccd", X"00000000", X"45ab17f8"),
		(X"429b0000", X"00000000", X"45ab88d1"),
		(X"429b3333", X"00000000", X"45abf9d0"),
		(X"429b6666", X"00000000", X"45ac6af4"),
		(X"429b999a", X"00000000", X"45acdc3e"),
		(X"429bcccd", X"00000000", X"45ad4dac"),
		(X"429c0000", X"00000000", X"45adbf40"),
		(X"429c3333", X"00000000", X"45ae30f9"),
		(X"429c6666", X"00000000", X"45aea2d7"),
		(X"429c999a", X"00000000", X"45af14da"),
		(X"429ccccd", X"00000000", X"45af8702"),
		(X"429d0000", X"00000000", X"45aff950"),
		(X"429d3333", X"00000000", X"45b06bc2"),
		(X"429d6666", X"00000000", X"45b0de5a"),
		(X"429d999a", X"00000000", X"45b15117"),
		(X"429dcccd", X"00000000", X"45b1c3f9"),
		(X"429e0000", X"00000000", X"45b23701"),
		(X"429e3333", X"00000000", X"45b2aa2d"),
		(X"429e6666", X"00000000", X"45b31d7f"),
		(X"429e999a", X"00000000", X"45b390f6"),
		(X"429ecccd", X"00000000", X"45b40492"),
		(X"429f0000", X"00000000", X"45b47853"),
		(X"429f3333", X"00000000", X"45b4ec39"),
		(X"429f6666", X"00000000", X"45b56045"),
		(X"429f999a", X"00000000", X"45b5d476"),
		(X"429fcccd", X"00000000", X"45b648cb"),
		(X"42a00000", X"00000000", X"45aa0553"),
		(X"42a03333", X"00000000", X"45aa71ce"),
		(X"42a06666", X"00000000", X"45aade6b"),
		(X"42a0999a", X"00000000", X"45ab4b2c"),
		(X"42a0cccd", X"00000000", X"45abb80e"),
		(X"42a10000", X"00000000", X"45ac2514"),
		(X"42a13333", X"00000000", X"45ac923c"),
		(X"42a16666", X"00000000", X"45acff86"),
		(X"42a1999a", X"00000000", X"45ad6cf3"),
		(X"42a1cccd", X"00000000", X"45adda83"),
		(X"42a20000", X"00000000", X"45ae4835"),
		(X"42a23333", X"00000000", X"45aeb60a"),
		(X"42a26666", X"00000000", X"45af2401"),
		(X"42a2999a", X"00000000", X"45af921b"),
		(X"42a2cccd", X"00000000", X"45b00057"),
		(X"42a30000", X"00000000", X"45b06eb6"),
		(X"42a33333", X"00000000", X"45b0dd38"),
		(X"42a36666", X"00000000", X"45b14bdc"),
		(X"42a3999a", X"00000000", X"45b1baa3"),
		(X"42a3cccd", X"00000000", X"45b2298c"),
		(X"42a40000", X"00000000", X"45b29898"),
		(X"42a43333", X"00000000", X"45b307c6"),
		(X"42a46666", X"00000000", X"45b37717"),
		(X"42a4999a", X"00000000", X"45b3e68a"),
		(X"42a4cccd", X"00000000", X"45b45620"),
		(X"42a50000", X"00000000", X"45b4c5d9"),
		(X"42a53333", X"00000000", X"45b535b4"),
		(X"42a56666", X"00000000", X"45b5a5b2"),
		(X"42a5999a", X"00000000", X"45b615d2"),
		(X"42a5cccd", X"00000000", X"45b68615"),
		(X"42a60000", X"00000000", X"45b6f67b"),
		(X"42a63333", X"00000000", X"45b76703"),
		(X"42a66666", X"00000000", X"45b7d7ad"),
		(X"42a6999a", X"00000000", X"45b8487a"),
		(X"42a6cccd", X"00000000", X"45b8b96a"),
		(X"42a70000", X"00000000", X"45b92a7c"),
		(X"42a73333", X"00000000", X"45b99bb1"),
		(X"42a76666", X"00000000", X"45ba0d09"),
		(X"42a7999a", X"00000000", X"45ba7e83"),
		(X"42a7cccd", X"00000000", X"45baf01f"),
		(X"42a80000", X"00000000", X"42927498"),
		(X"42a83333", X"00000000", X"4292b449"),
		(X"42a86666", X"00000000", X"4292f406"),
		(X"42a8999a", X"00000000", X"429333ce"),
		(X"42a8cccd", X"00000000", X"429373a1"),
		(X"42a90000", X"00000000", X"4293b381"),
		(X"42a93333", X"00000000", X"4293f36b"),
		(X"42a96666", X"00000000", X"42943362"),
		(X"42a9999a", X"00000000", X"42947364"),
		(X"42a9cccd", X"00000000", X"4294b372"),
		(X"42aa0000", X"00000000", X"4294f38b"),
		(X"42aa3333", X"00000000", X"429533b0"),
		(X"42aa6666", X"00000000", X"429573e0"),
		(X"42aa999a", X"00000000", X"4295b41c"),
		(X"42aacccd", X"00000000", X"4295f464"),
		(X"42ab0000", X"00000000", X"429634b7"),
		(X"42ab3333", X"00000000", X"42967516"),
		(X"42ab6666", X"00000000", X"4296b580"),
		(X"42ab999a", X"00000000", X"4296f5f6"),
		(X"42abcccd", X"00000000", X"42973678"),
		(X"42ac0000", X"00000000", X"42977705"),
		(X"42ac3333", X"00000000", X"4297b79e"),
		(X"42ac6666", X"00000000", X"4297f843"),
		(X"42ac999a", X"00000000", X"429838f3"),
		(X"42accccd", X"00000000", X"429879ae"),
		(X"42ad0000", X"00000000", X"4298ba76"),
		(X"42ad3333", X"00000000", X"4298fb49"),
		(X"42ad6666", X"00000000", X"42993c27"),
		(X"42ad999a", X"00000000", X"42997d11"),
		(X"42adcccd", X"00000000", X"4299be07"),
		(X"42ae0000", X"00000000", X"4299ff08"),
		(X"42ae3333", X"00000000", X"429a4015"),
		(X"42ae6666", X"00000000", X"429a812d"),
		(X"42ae999a", X"00000000", X"429ac251"),
		(X"42aecccd", X"00000000", X"429b0381"),
		(X"42af0000", X"00000000", X"429b44bc"),
		(X"42af3333", X"00000000", X"429b8603"),
		(X"42af6666", X"00000000", X"429bc756"),
		(X"42af999a", X"00000000", X"429c08b4"),
		(X"42afcccd", X"00000000", X"429c4a1e"),
		(X"42b00000", X"00000000", X"c5c9ae29"),
		(X"42b03333", X"00000000", X"c5ca23f8"),
		(X"42b06666", X"00000000", X"c5ca99e9"),
		(X"42b0999a", X"00000000", X"c5cb0ffd"),
		(X"42b0cccd", X"00000000", X"c5cb8633"),
		(X"42b10000", X"00000000", X"c5cbfc8b"),
		(X"42b13333", X"00000000", X"c5cc7306"),
		(X"42b16666", X"00000000", X"c5cce9a3"),
		(X"42b1999a", X"00000000", X"c5cd6063"),
		(X"42b1cccd", X"00000000", X"c5cdd745"),
		(X"42b20000", X"00000000", X"c5ce4e49"),
		(X"42b23333", X"00000000", X"c5cec570"),
		(X"42b26666", X"00000000", X"c5cf3cb9"),
		(X"42b2999a", X"00000000", X"c5cfb424"),
		(X"42b2cccd", X"00000000", X"c5d02bb2"),
		(X"42b30000", X"00000000", X"c5d0a362"),
		(X"42b33333", X"00000000", X"c5d11b34"),
		(X"42b36666", X"00000000", X"c5d19329"),
		(X"42b3999a", X"00000000", X"c5d20b40"),
		(X"42b3cccd", X"00000000", X"c5d2837a"),
		(X"42b40000", X"00000000", X"c5d2fbd6"),
		(X"42b43333", X"00000000", X"c5d37454"),
		(X"42b46666", X"00000000", X"c5d3ecf5"),
		(X"42b4999a", X"00000000", X"c5d465b8"),
		(X"42b4cccd", X"00000000", X"c5d4de9d"),
		(X"42b50000", X"00000000", X"c5d557a5"),
		(X"42b53333", X"00000000", X"c5d5d0cf"),
		(X"42b56666", X"00000000", X"c5d64a1c"),
		(X"42b5999a", X"00000000", X"c5d6c38b"),
		(X"42b5cccd", X"00000000", X"c5d73d1c"),
		(X"42b60000", X"00000000", X"c5d7b6d0"),
		(X"42b63333", X"00000000", X"c5d830a6"),
		(X"42b66666", X"00000000", X"c5d8aa9e"),
		(X"42b6999a", X"00000000", X"c5d924b9"),
		(X"42b6cccd", X"00000000", X"c5d99ef6"),
		(X"42b70000", X"00000000", X"c5da1955"),
		(X"42b73333", X"00000000", X"c5da93d7"),
		(X"42b76666", X"00000000", X"c5db0e7b"),
		(X"42b7999a", X"00000000", X"c5db8942"),
		(X"42b7cccd", X"00000000", X"c5dc042b"),
		(X"42b80000", X"00000000", X"c5ef8e74"),
		(X"42b83333", X"00000000", X"c5f0143e"),
		(X"42b86666", X"00000000", X"c5f09a2e"),
		(X"42b8999a", X"00000000", X"c5f12043"),
		(X"42b8cccd", X"00000000", X"c5f1a67e"),
		(X"42b90000", X"00000000", X"c5f22cde"),
		(X"42b93333", X"00000000", X"c5f2b363"),
		(X"42b96666", X"00000000", X"c5f33a0d"),
		(X"42b9999a", X"00000000", X"c5f3c0dd"),
		(X"42b9cccd", X"00000000", X"c5f447d2"),
		(X"42ba0000", X"00000000", X"c5f4ceed"),
		(X"42ba3333", X"00000000", X"c5f5562d"),
		(X"42ba6666", X"00000000", X"c5f5dd92"),
		(X"42ba999a", X"00000000", X"c5f6651c"),
		(X"42bacccd", X"00000000", X"c5f6eccc"),
		(X"42bb0000", X"00000000", X"c5f774a1"),
		(X"42bb3333", X"00000000", X"c5f7fc9b"),
		(X"42bb6666", X"00000000", X"c5f884bb"),
		(X"42bb999a", X"00000000", X"c5f90d00"),
		(X"42bbcccd", X"00000000", X"c5f9956a"),
		(X"42bc0000", X"00000000", X"c5fa1dfa"),
		(X"42bc3333", X"00000000", X"c5faa6af"),
		(X"42bc6666", X"00000000", X"c5fb2f89"),
		(X"42bc999a", X"00000000", X"c5fbb889"),
		(X"42bccccd", X"00000000", X"c5fc41ae"),
		(X"42bd0000", X"00000000", X"c5fccaf8"),
		(X"42bd3333", X"00000000", X"c5fd5467"),
		(X"42bd6666", X"00000000", X"c5fdddfc"),
		(X"42bd999a", X"00000000", X"c5fe67b6"),
		(X"42bdcccd", X"00000000", X"c5fef196"),
		(X"42be0000", X"00000000", X"c5ff7b9b"),
		(X"42be3333", X"00000000", X"c60002e3"),
		(X"42be6666", X"00000000", X"c600480a"),
		(X"42be999a", X"00000000", X"c6008d45"),
		(X"42becccd", X"00000000", X"c600d292"),
		(X"42bf0000", X"00000000", X"c60117f1"),
		(X"42bf3333", X"00000000", X"c6015d64"),
		(X"42bf6666", X"00000000", X"c601a2e9"),
		(X"42bf999a", X"00000000", X"c601e881"),
		(X"42bfcccd", X"00000000", X"c6022e2b"),
		(X"42c00000", X"00000000", X"c4a19db5"),
		(X"42c03333", X"00000000", X"c4a1f58c"),
		(X"42c06666", X"00000000", X"c4a24d7c"),
		(X"42c0999a", X"00000000", X"c4a2a583"),
		(X"42c0cccd", X"00000000", X"c4a2fda2"),
		(X"42c10000", X"00000000", X"c4a355d9"),
		(X"42c13333", X"00000000", X"c4a3ae27"),
		(X"42c16666", X"00000000", X"c4a4068e"),
		(X"42c1999a", X"00000000", X"c4a45f0c"),
		(X"42c1cccd", X"00000000", X"c4a4b7a2"),
		(X"42c20000", X"00000000", X"c4a51050"),
		(X"42c23333", X"00000000", X"c4a56916"),
		(X"42c26666", X"00000000", X"c4a5c1f4"),
		(X"42c2999a", X"00000000", X"c4a61aea"),
		(X"42c2cccd", X"00000000", X"c4a673f7"),
		(X"42c30000", X"00000000", X"c4a6cd1c"),
		(X"42c33333", X"00000000", X"c4a72659"),
		(X"42c36666", X"00000000", X"c4a77fae"),
		(X"42c3999a", X"00000000", X"c4a7d91b"),
		(X"42c3cccd", X"00000000", X"c4a832a0"),
		(X"42c40000", X"00000000", X"c4a88c3c"),
		(X"42c43333", X"00000000", X"c4a8e5f0"),
		(X"42c46666", X"00000000", X"c4a93fbc"),
		(X"42c4999a", X"00000000", X"c4a999a0"),
		(X"42c4cccd", X"00000000", X"c4a9f39c"),
		(X"42c50000", X"00000000", X"c4aa4db0"),
		(X"42c53333", X"00000000", X"c4aaa7db"),
		(X"42c56666", X"00000000", X"c4ab021f"),
		(X"42c5999a", X"00000000", X"c4ab5c7a"),
		(X"42c5cccd", X"00000000", X"c4abb6ed"),
		(X"42c60000", X"00000000", X"c4ac1177"),
		(X"42c63333", X"00000000", X"c4ac6c1a"),
		(X"42c66666", X"00000000", X"c4acc6d5"),
		(X"42c6999a", X"00000000", X"c4ad21a7"),
		(X"42c6cccd", X"00000000", X"c4ad7c91"),
		(X"42c70000", X"00000000", X"c4add793"),
		(X"42c73333", X"00000000", X"c4ae32ad"),
		(X"42c76666", X"00000000", X"c4ae8ddf"),
		(X"42c7999a", X"00000000", X"c4aee928"),
		(X"42c7cccd", X"00000000", X"c4af448a"),
		(X"42c80000", X"00000000", X"45ed282e"),
		(X"42c83333", X"00000000", X"45eda144"),
		(X"42c86666", X"00000000", X"45ee1a78"),
		(X"42c8999a", X"00000000", X"45ee93cc"),
		(X"42c8cccd", X"00000000", X"45ef0d3e"),
		(X"42c90000", X"00000000", X"45ef86cf"),
		(X"42c93333", X"00000000", X"45f0007f"),
		(X"42c96666", X"00000000", X"45f07a4e"),
		(X"42c9999a", X"00000000", X"45f0f43c"),
		(X"42c9cccd", X"00000000", X"45f16e49"),
		(X"42ca0000", X"00000000", X"45f1e875"),
		(X"42ca3333", X"00000000", X"45f262bf"),
		(X"42ca6666", X"00000000", X"45f2dd28"),
		(X"42ca999a", X"00000000", X"45f357b1"),
		(X"42cacccd", X"00000000", X"45f3d258"),
		(X"42cb0000", X"00000000", X"45f44d1e"),
		(X"42cb3333", X"00000000", X"45f4c803"),
		(X"42cb6666", X"00000000", X"45f54306"),
		(X"42cb999a", X"00000000", X"45f5be29"),
		(X"42cbcccd", X"00000000", X"45f6396a"),
		(X"42cc0000", X"00000000", X"45f6b4cb"),
		(X"42cc3333", X"00000000", X"45f7304a"),
		(X"42cc6666", X"00000000", X"45f7abe8"),
		(X"42cc999a", X"00000000", X"45f827a5"),
		(X"42cccccd", X"00000000", X"45f8a381"),
		(X"42cd0000", X"00000000", X"45f91f7c"),
		(X"42cd3333", X"00000000", X"45f99b96"),
		(X"42cd6666", X"00000000", X"45fa17ce"),
		(X"42cd999a", X"00000000", X"45fa9426"),
		(X"42cdcccd", X"00000000", X"45fb109c"),
		(X"42ce0000", X"00000000", X"45fb8d31"),
		(X"42ce3333", X"00000000", X"45fc09e5"),
		(X"42ce6666", X"00000000", X"45fc86b8"),
		(X"42ce999a", X"00000000", X"45fd03aa"),
		(X"42cecccd", X"00000000", X"45fd80bb"),
		(X"42cf0000", X"00000000", X"45fdfdea"),
		(X"42cf3333", X"00000000", X"45fe7b39"),
		(X"42cf6666", X"00000000", X"45fef8a6"),
		(X"42cf999a", X"00000000", X"45ff7632"),
		(X"42cfcccd", X"00000000", X"45fff3de"),
		(X"42d00000", X"00000000", X"462314cf"),
		(X"42d03333", X"00000000", X"462364ef"),
		(X"42d06666", X"00000000", X"4623b522"),
		(X"42d0999a", X"00000000", X"46240569"),
		(X"42d0cccd", X"00000000", X"462455c4"),
		(X"42d10000", X"00000000", X"4624a633"),
		(X"42d13333", X"00000000", X"4624f6b5"),
		(X"42d16666", X"00000000", X"4625474b"),
		(X"42d1999a", X"00000000", X"462597f4"),
		(X"42d1cccd", X"00000000", X"4625e8b2"),
		(X"42d20000", X"00000000", X"46263982"),
		(X"42d23333", X"00000000", X"46268a67"),
		(X"42d26666", X"00000000", X"4626db5f"),
		(X"42d2999a", X"00000000", X"46272c6b"),
		(X"42d2cccd", X"00000000", X"46277d8b"),
		(X"42d30000", X"00000000", X"4627cebe"),
		(X"42d33333", X"00000000", X"46282005"),
		(X"42d36666", X"00000000", X"4628715f"),
		(X"42d3999a", X"00000000", X"4628c2cd"),
		(X"42d3cccd", X"00000000", X"4629144f"),
		(X"42d40000", X"00000000", X"462965e5"),
		(X"42d43333", X"00000000", X"4629b78e"),
		(X"42d46666", X"00000000", X"462a094b"),
		(X"42d4999a", X"00000000", X"462a5b1b"),
		(X"42d4cccd", X"00000000", X"462aacff"),
		(X"42d50000", X"00000000", X"462afef7"),
		(X"42d53333", X"00000000", X"462b5103"),
		(X"42d56666", X"00000000", X"462ba322"),
		(X"42d5999a", X"00000000", X"462bf555"),
		(X"42d5cccd", X"00000000", X"462c479b"),
		(X"42d60000", X"00000000", X"462c99f5"),
		(X"42d63333", X"00000000", X"462cec63"),
		(X"42d66666", X"00000000", X"462d3ee5"),
		(X"42d6999a", X"00000000", X"462d917a"),
		(X"42d6cccd", X"00000000", X"462de423"),
		(X"42d70000", X"00000000", X"462e36df"),
		(X"42d73333", X"00000000", X"462e89af"),
		(X"42d76666", X"00000000", X"462edc93"),
		(X"42d7999a", X"00000000", X"462f2f8b"),
		(X"42d7cccd", X"00000000", X"462f8296"),
		(X"42d80000", X"00000000", X"45522a2c"),
		(X"42d83333", X"00000000", X"45528d0d"),
		(X"42d86666", X"00000000", X"4552f005"),
		(X"42d8999a", X"00000000", X"45535315"),
		(X"42d8cccd", X"00000000", X"4553b63c"),
		(X"42d90000", X"00000000", X"45541979"),
		(X"42d93333", X"00000000", X"45547ccf"),
		(X"42d96666", X"00000000", X"4554e03b"),
		(X"42d9999a", X"00000000", X"455543bf"),
		(X"42d9cccd", X"00000000", X"4555a75a"),
		(X"42da0000", X"00000000", X"45560b0c"),
		(X"42da3333", X"00000000", X"45566ed5"),
		(X"42da6666", X"00000000", X"4556d2b6"),
		(X"42da999a", X"00000000", X"455736ae"),
		(X"42dacccd", X"00000000", X"45579abd"),
		(X"42db0000", X"00000000", X"4557fee3"),
		(X"42db3333", X"00000000", X"45586321"),
		(X"42db6666", X"00000000", X"4558c776"),
		(X"42db999a", X"00000000", X"45592be2"),
		(X"42dbcccd", X"00000000", X"45599065"),
		(X"42dc0000", X"00000000", X"4559f500"),
		(X"42dc3333", X"00000000", X"455a59b2"),
		(X"42dc6666", X"00000000", X"455abe7b"),
		(X"42dc999a", X"00000000", X"455b235b"),
		(X"42dccccd", X"00000000", X"455b8852"),
		(X"42dd0000", X"00000000", X"455bed61"),
		(X"42dd3333", X"00000000", X"455c5287"),
		(X"42dd6666", X"00000000", X"455cb7c4"),
		(X"42dd999a", X"00000000", X"455d1d19"),
		(X"42ddcccd", X"00000000", X"455d8284"),
		(X"42de0000", X"00000000", X"455de807"),
		(X"42de3333", X"00000000", X"455e4da1"),
		(X"42de6666", X"00000000", X"455eb353"),
		(X"42de999a", X"00000000", X"455f191c"),
		(X"42decccd", X"00000000", X"455f7efb"),
		(X"42df0000", X"00000000", X"455fe4f3"),
		(X"42df3333", X"00000000", X"45604b01"),
		(X"42df6666", X"00000000", X"4560b126"),
		(X"42df999a", X"00000000", X"45611763"),
		(X"42dfcccd", X"00000000", X"45617db7"),
		(X"42e00000", X"00000000", X"c5fe7a72"),
		(X"42e03333", X"00000000", X"c5feef3b"),
		(X"42e06666", X"00000000", X"c5ff641f"),
		(X"42e0999a", X"00000000", X"c5ffd91d"),
		(X"42e0cccd", X"00000000", X"c600271b"),
		(X"42e10000", X"00000000", X"c60061b5"),
		(X"42e13333", X"00000000", X"c6009c5d"),
		(X"42e16666", X"00000000", X"c600d712"),
		(X"42e1999a", X"00000000", X"c60111d4"),
		(X"42e1cccd", X"00000000", X"c6014ca3"),
		(X"42e20000", X"00000000", X"c6018780"),
		(X"42e23333", X"00000000", X"c601c26b"),
		(X"42e26666", X"00000000", X"c601fd63"),
		(X"42e2999a", X"00000000", X"c6023868"),
		(X"42e2cccd", X"00000000", X"c602737a"),
		(X"42e30000", X"00000000", X"c602ae9a"),
		(X"42e33333", X"00000000", X"c602e9c7"),
		(X"42e36666", X"00000000", X"c6032502"),
		(X"42e3999a", X"00000000", X"c603604a"),
		(X"42e3cccd", X"00000000", X"c6039ba0"),
		(X"42e40000", X"00000000", X"c603d703"),
		(X"42e43333", X"00000000", X"c6041273"),
		(X"42e46666", X"00000000", X"c6044df0"),
		(X"42e4999a", X"00000000", X"c604897b"),
		(X"42e4cccd", X"00000000", X"c604c514"),
		(X"42e50000", X"00000000", X"c60500ba"),
		(X"42e53333", X"00000000", X"c6053c6d"),
		(X"42e56666", X"00000000", X"c605782d"),
		(X"42e5999a", X"00000000", X"c605b3fb"),
		(X"42e5cccd", X"00000000", X"c605efd7"),
		(X"42e60000", X"00000000", X"c6062bbf"),
		(X"42e63333", X"00000000", X"c60667b5"),
		(X"42e66666", X"00000000", X"c606a3b9"),
		(X"42e6999a", X"00000000", X"c606dfca"),
		(X"42e6cccd", X"00000000", X"c6071be8"),
		(X"42e70000", X"00000000", X"c6075814"),
		(X"42e73333", X"00000000", X"c607944d"),
		(X"42e76666", X"00000000", X"c607d093"),
		(X"42e7999a", X"00000000", X"c6080ce7"),
		(X"42e7cccd", X"00000000", X"c6084948"),
		(X"42e80000", X"00000000", X"c64f3d5b"),
		(X"42e83333", X"00000000", X"c64f9911"),
		(X"42e86666", X"00000000", X"c64ff4db"),
		(X"42e8999a", X"00000000", X"c65050ba"),
		(X"42e8cccd", X"00000000", X"c650acad"),
		(X"42e90000", X"00000000", X"c65108b4"),
		(X"42e93333", X"00000000", X"c65164cf"),
		(X"42e96666", X"00000000", X"c651c0ff"),
		(X"42e9999a", X"00000000", X"c6521d43"),
		(X"42e9cccd", X"00000000", X"c652799b"),
		(X"42ea0000", X"00000000", X"c652d607"),
		(X"42ea3333", X"00000000", X"c6533288"),
		(X"42ea6666", X"00000000", X"c6538f1d"),
		(X"42ea999a", X"00000000", X"c653ebc7"),
		(X"42eacccd", X"00000000", X"c6544884"),
		(X"42eb0000", X"00000000", X"c654a556"),
		(X"42eb3333", X"00000000", X"c655023c"),
		(X"42eb6666", X"00000000", X"c6555f36"),
		(X"42eb999a", X"00000000", X"c655bc45"),
		(X"42ebcccd", X"00000000", X"c6561968"),
		(X"42ec0000", X"00000000", X"c656769f"),
		(X"42ec3333", X"00000000", X"c656d3eb"),
		(X"42ec6666", X"00000000", X"c657314b"),
		(X"42ec999a", X"00000000", X"c6578ebf"),
		(X"42eccccd", X"00000000", X"c657ec47"),
		(X"42ed0000", X"00000000", X"c65849e3"),
		(X"42ed3333", X"00000000", X"c658a794"),
		(X"42ed6666", X"00000000", X"c6590559"),
		(X"42ed999a", X"00000000", X"c6596333"),
		(X"42edcccd", X"00000000", X"c659c121"),
		(X"42ee0000", X"00000000", X"c65a1f23"),
		(X"42ee3333", X"00000000", X"c65a7d39"),
		(X"42ee6666", X"00000000", X"c65adb63"),
		(X"42ee999a", X"00000000", X"c65b39a2"),
		(X"42eecccd", X"00000000", X"c65b97f5"),
		(X"42ef0000", X"00000000", X"c65bf65d"),
		(X"42ef3333", X"00000000", X"c65c54d8"),
		(X"42ef6666", X"00000000", X"c65cb368"),
		(X"42ef999a", X"00000000", X"c65d120c"),
		(X"42efcccd", X"00000000", X"c65d70c5"),
		(X"42f00000", X"00000000", X"c5b9641e"),
		(X"42f03333", X"00000000", X"c5b9b3a6"),
		(X"42f06666", X"00000000", X"c5ba0340"),
		(X"42f0999a", X"00000000", X"c5ba52ea"),
		(X"42f0cccd", X"00000000", X"c5baa2a6"),
		(X"42f10000", X"00000000", X"c5baf273"),
		(X"42f13333", X"00000000", X"c5bb4251"),
		(X"42f16666", X"00000000", X"c5bb9240"),
		(X"42f1999a", X"00000000", X"c5bbe23f"),
		(X"42f1cccd", X"00000000", X"c5bc3250"),
		(X"42f20000", X"00000000", X"c5bc8272"),
		(X"42f23333", X"00000000", X"c5bcd2a5"),
		(X"42f26666", X"00000000", X"c5bd22e9"),
		(X"42f2999a", X"00000000", X"c5bd733f"),
		(X"42f2cccd", X"00000000", X"c5bdc3a5"),
		(X"42f30000", X"00000000", X"c5be141c"),
		(X"42f33333", X"00000000", X"c5be64a4"),
		(X"42f36666", X"00000000", X"c5beb53d"),
		(X"42f3999a", X"00000000", X"c5bf05e8"),
		(X"42f3cccd", X"00000000", X"c5bf56a3"),
		(X"42f40000", X"00000000", X"c5bfa770"),
		(X"42f43333", X"00000000", X"c5bff84d"),
		(X"42f46666", X"00000000", X"c5c0493c"),
		(X"42f4999a", X"00000000", X"c5c09a3b"),
		(X"42f4cccd", X"00000000", X"c5c0eb4c"),
		(X"42f50000", X"00000000", X"c5c13c6d"),
		(X"42f53333", X"00000000", X"c5c18da0"),
		(X"42f56666", X"00000000", X"c5c1dee4"),
		(X"42f5999a", X"00000000", X"c5c23039"),
		(X"42f5cccd", X"00000000", X"c5c2819f"),
		(X"42f60000", X"00000000", X"c5c2d315"),
		(X"42f63333", X"00000000", X"c5c3249d"),
		(X"42f66666", X"00000000", X"c5c37636"),
		(X"42f6999a", X"00000000", X"c5c3c7e0"),
		(X"42f6cccd", X"00000000", X"c5c4199b"),
		(X"42f70000", X"00000000", X"c5c46b68"),
		(X"42f73333", X"00000000", X"c5c4bd45"),
		(X"42f76666", X"00000000", X"c5c50f33"),
		(X"42f7999a", X"00000000", X"c5c56132"),
		(X"42f7cccd", X"00000000", X"c5c5b343"),
		(X"42f80000", X"00000000", X"4602c6c1"),
		(X"42f83333", X"00000000", X"4602fc93"),
		(X"42f86666", X"00000000", X"4603326f"),
		(X"42f8999a", X"00000000", X"46036857"),
		(X"42f8cccd", X"00000000", X"46039e4a"),
		(X"42f90000", X"00000000", X"4603d449"),
		(X"42f93333", X"00000000", X"46040a52"),
		(X"42f96666", X"00000000", X"46044066"),
		(X"42f9999a", X"00000000", X"46047685"),
		(X"42f9cccd", X"00000000", X"4604acaf"),
		(X"42fa0000", X"00000000", X"4604e2e5"),
		(X"42fa3333", X"00000000", X"46051925"),
		(X"42fa6666", X"00000000", X"46054f71"),
		(X"42fa999a", X"00000000", X"460585c8"),
		(X"42facccd", X"00000000", X"4605bc29"),
		(X"42fb0000", X"00000000", X"4605f296"),
		(X"42fb3333", X"00000000", X"4606290e"),
		(X"42fb6666", X"00000000", X"46065f91"),
		(X"42fb999a", X"00000000", X"4606961e"),
		(X"42fbcccd", X"00000000", X"4606ccb7"),
		(X"42fc0000", X"00000000", X"4607035c"),
		(X"42fc3333", X"00000000", X"46073a0b"),
		(X"42fc6666", X"00000000", X"460770c5"),
		(X"42fc999a", X"00000000", X"4607a78a"),
		(X"42fccccd", X"00000000", X"4607de5a"),
		(X"42fd0000", X"00000000", X"46081536"),
		(X"42fd3333", X"00000000", X"46084c1c"),
		(X"42fd6666", X"00000000", X"4608830e"),
		(X"42fd999a", X"00000000", X"4608ba0a"),
		(X"42fdcccd", X"00000000", X"4608f112"),
		(X"42fe0000", X"00000000", X"46092825"),
		(X"42fe3333", X"00000000", X"46095f43"),
		(X"42fe6666", X"00000000", X"4609966b"),
		(X"42fe999a", X"00000000", X"4609cd9f"),
		(X"42fecccd", X"00000000", X"460a04de"),
		(X"42ff0000", X"00000000", X"460a3c28"),
		(X"42ff3333", X"00000000", X"460a737d"),
		(X"42ff6666", X"00000000", X"460aaade"),
		(X"42ff999a", X"00000000", X"460ae249"),
		(X"42ffcccd", X"00000000", X"460b19bf"),
		(X"43000000", X"00000000", X"46808000"),
		(X"4300199a", X"00000000", X"4680b352"),
		(X"43003333", X"00000000", X"4680e6ae"),
		(X"43004ccd", X"00000000", X"46811a14"),
		(X"43006666", X"00000000", X"46814d85"),
		(X"43008000", X"00000000", X"46818100"),
		(X"4300999a", X"00000000", X"4681b485"),
		(X"4300b333", X"00000000", X"4681e814"),
		(X"4300cccd", X"00000000", X"46821bae"),
		(X"4300e666", X"00000000", X"46824f52"),
		(X"43010000", X"00000000", X"46828300"),
		(X"4301199a", X"00000000", X"4682b6b8"),
		(X"43013333", X"00000000", X"4682ea7b"),
		(X"43014ccd", X"00000000", X"46831e48"),
		(X"43016666", X"00000000", X"4683521f"),
		(X"43018000", X"00000000", X"46838600"),
		(X"4301999a", X"00000000", X"4683b9ec"),
		(X"4301b333", X"00000000", X"4683ede1"),
		(X"4301cccd", X"00000000", X"468421e1"),
		(X"4301e666", X"00000000", X"468455ec"),
		(X"43020000", X"00000000", X"46848a00"),
		(X"4302199a", X"00000000", X"4684be1f"),
		(X"43023333", X"00000000", X"4684f248"),
		(X"43024ccd", X"00000000", X"4685267b"),
		(X"43026666", X"00000000", X"46855ab8"),
		(X"43028000", X"00000000", X"46858f00"),
		(X"4302999a", X"00000000", X"4685c352"),
		(X"4302b333", X"00000000", X"4685f7ae"),
		(X"4302cccd", X"00000000", X"46862c14"),
		(X"4302e666", X"00000000", X"46866085"),
		(X"43030000", X"00000000", X"46869500"),
		(X"4303199a", X"00000000", X"4686c985"),
		(X"43033333", X"00000000", X"4686fe14"),
		(X"43034ccd", X"00000000", X"468732ae"),
		(X"43036666", X"00000000", X"46876752"),
		(X"43038000", X"00000000", X"46879c00"),
		(X"4303999a", X"00000000", X"4687d0b8"),
		(X"4303b333", X"00000000", X"4688057b"),
		(X"4303cccd", X"00000000", X"46883a48"),
		(X"4303e666", X"00000000", X"46886f1f"),
		(X"43040000", X"00000000", X"461420e9"),
		(X"4304199a", X"00000000", X"46145a30"),
		(X"43043333", X"00000000", X"46149382"),
		(X"43044ccd", X"00000000", X"4614ccdf"),
		(X"43046666", X"00000000", X"46150647"),
		(X"43048000", X"00000000", X"46153fbb"),
		(X"4304999a", X"00000000", X"46157939"),
		(X"4304b333", X"00000000", X"4615b2c3"),
		(X"4304cccd", X"00000000", X"4615ec57"),
		(X"4304e666", X"00000000", X"461625f7"),
		(X"43050000", X"00000000", X"46165fa1"),
		(X"4305199a", X"00000000", X"46169957"),
		(X"43053333", X"00000000", X"4616d318"),
		(X"43054ccd", X"00000000", X"46170ce4"),
		(X"43056666", X"00000000", X"461746ba"),
		(X"43058000", X"00000000", X"4617809c"),
		(X"4305999a", X"00000000", X"4617ba89"),
		(X"4305b333", X"00000000", X"4617f482"),
		(X"4305cccd", X"00000000", X"46182e85"),
		(X"4305e666", X"00000000", X"46186893"),
		(X"43060000", X"00000000", X"4618a2ac"),
		(X"4306199a", X"00000000", X"4618dcd1"),
		(X"43063333", X"00000000", X"46191700"),
		(X"43064ccd", X"00000000", X"4619513b"),
		(X"43066666", X"00000000", X"46198b80"),
		(X"43068000", X"00000000", X"4619c5d1"),
		(X"4306999a", X"00000000", X"461a002c"),
		(X"4306b333", X"00000000", X"461a3a93"),
		(X"4306cccd", X"00000000", X"461a7505"),
		(X"4306e666", X"00000000", X"461aaf82"),
		(X"43070000", X"00000000", X"461aea0a"),
		(X"4307199a", X"00000000", X"461b249d"),
		(X"43073333", X"00000000", X"461b5f3b"),
		(X"43074ccd", X"00000000", X"461b99e4"),
		(X"43076666", X"00000000", X"461bd498"),
		(X"43078000", X"00000000", X"461c0f57"),
		(X"4307999a", X"00000000", X"461c4a22"),
		(X"4307b333", X"00000000", X"461c84f7"),
		(X"4307cccd", X"00000000", X"461cbfd8"),
		(X"4307e666", X"00000000", X"461cfac3"),
		(X"43080000", X"00000000", X"c5ee686a"),
		(X"4308199a", X"00000000", X"c5eec29a"),
		(X"43083333", X"00000000", X"c5ef1cdb"),
		(X"43084ccd", X"00000000", X"c5ef772d"),
		(X"43086666", X"00000000", X"c5efd190"),
		(X"43088000", X"00000000", X"c5f02c04"),
		(X"4308999a", X"00000000", X"c5f08689"),
		(X"4308b333", X"00000000", X"c5f0e11f"),
		(X"4308cccd", X"00000000", X"c5f13bc6"),
		(X"4308e666", X"00000000", X"c5f1967e"),
		(X"43090000", X"00000000", X"c5f1f148"),
		(X"4309199a", X"00000000", X"c5f24c22"),
		(X"43093333", X"00000000", X"c5f2a70d"),
		(X"43094ccd", X"00000000", X"c5f3020a"),
		(X"43096666", X"00000000", X"c5f35d17"),
		(X"43098000", X"00000000", X"c5f3b836"),
		(X"4309999a", X"00000000", X"c5f41365"),
		(X"4309b333", X"00000000", X"c5f46ea6"),
		(X"4309cccd", X"00000000", X"c5f4c9f7"),
		(X"4309e666", X"00000000", X"c5f5255a"),
		(X"430a0000", X"00000000", X"c5f580ce"),
		(X"430a199a", X"00000000", X"c5f5dc52"),
		(X"430a3333", X"00000000", X"c5f637e8"),
		(X"430a4ccd", X"00000000", X"c5f6938f"),
		(X"430a6666", X"00000000", X"c5f6ef47"),
		(X"430a8000", X"00000000", X"c5f74b10"),
		(X"430a999a", X"00000000", X"c5f7a6ea"),
		(X"430ab333", X"00000000", X"c5f802d5"),
		(X"430acccd", X"00000000", X"c5f85ed1"),
		(X"430ae666", X"00000000", X"c5f8bade"),
		(X"430b0000", X"00000000", X"c5f916fc"),
		(X"430b199a", X"00000000", X"c5f9732b"),
		(X"430b3333", X"00000000", X"c5f9cf6b"),
		(X"430b4ccd", X"00000000", X"c5fa2bbd"),
		(X"430b6666", X"00000000", X"c5fa881f"),
		(X"430b8000", X"00000000", X"c5fae492"),
		(X"430b999a", X"00000000", X"c5fb4117"),
		(X"430bb333", X"00000000", X"c5fb9dac"),
		(X"430bcccd", X"00000000", X"c5fbfa53"),
		(X"430be666", X"00000000", X"c5fc570a"),
		(X"430c0000", X"00000000", X"c6970bb5"),
		(X"430c199a", X"00000000", X"c6974311"),
		(X"430c3333", X"00000000", X"c6977a77"),
		(X"430c4ccd", X"00000000", X"c697b1e7"),
		(X"430c6666", X"00000000", X"c697e962"),
		(X"430c8000", X"00000000", X"c69820e6"),
		(X"430c999a", X"00000000", X"c6985875"),
		(X"430cb333", X"00000000", X"c698900e"),
		(X"430ccccd", X"00000000", X"c698c7b1"),
		(X"430ce666", X"00000000", X"c698ff5e"),
		(X"430d0000", X"00000000", X"c6993715"),
		(X"430d199a", X"00000000", X"c6996ed6"),
		(X"430d3333", X"00000000", X"c699a6a2"),
		(X"430d4ccd", X"00000000", X"c699de77"),
		(X"430d6666", X"00000000", X"c69a1657"),
		(X"430d8000", X"00000000", X"c69a4e41"),
		(X"430d999a", X"00000000", X"c69a8635"),
		(X"430db333", X"00000000", X"c69abe33"),
		(X"430dcccd", X"00000000", X"c69af63c"),
		(X"430de666", X"00000000", X"c69b2e4e"),
		(X"430e0000", X"00000000", X"c69b666b"),
		(X"430e199a", X"00000000", X"c69b9e92"),
		(X"430e3333", X"00000000", X"c69bd6c2"),
		(X"430e4ccd", X"00000000", X"c69c0efe"),
		(X"430e6666", X"00000000", X"c69c4743"),
		(X"430e8000", X"00000000", X"c69c7f92"),
		(X"430e999a", X"00000000", X"c69cb7eb"),
		(X"430eb333", X"00000000", X"c69cf04f"),
		(X"430ecccd", X"00000000", X"c69d28bd"),
		(X"430ee666", X"00000000", X"c69d6135"),
		(X"430f0000", X"00000000", X"c69d99b7"),
		(X"430f199a", X"00000000", X"c69dd243"),
		(X"430f3333", X"00000000", X"c69e0ad9"),
		(X"430f4ccd", X"00000000", X"c69e4379"),
		(X"430f6666", X"00000000", X"c69e7c24"),
		(X"430f8000", X"00000000", X"c69eb4d9"),
		(X"430f999a", X"00000000", X"c69eed97"),
		(X"430fb333", X"00000000", X"c69f2660"),
		(X"430fcccd", X"00000000", X"c69f5f33"),
		(X"430fe666", X"00000000", X"c69f9811"),
		(X"43100000", X"00000000", X"c652a7d1"),
		(X"4310199a", X"00000000", X"c652f2f1"),
		(X"43103333", X"00000000", X"c6533e1f"),
		(X"43104ccd", X"00000000", X"c653895a"),
		(X"43106666", X"00000000", X"c653d4a2"),
		(X"43108000", X"00000000", X"c6541ff8"),
		(X"4310999a", X"00000000", X"c6546b5b"),
		(X"4310b333", X"00000000", X"c654b6cc"),
		(X"4310cccd", X"00000000", X"c655024a"),
		(X"4310e666", X"00000000", X"c6554dd5"),
		(X"43110000", X"00000000", X"c655996e"),
		(X"4311199a", X"00000000", X"c655e514"),
		(X"43113333", X"00000000", X"c65630c7"),
		(X"43114ccd", X"00000000", X"c6567c88"),
		(X"43116666", X"00000000", X"c656c856"),
		(X"43118000", X"00000000", X"c6571432"),
		(X"4311999a", X"00000000", X"c657601b"),
		(X"4311b333", X"00000000", X"c657ac11"),
		(X"4311cccd", X"00000000", X"c657f815"),
		(X"4311e666", X"00000000", X"c6584426"),
		(X"43120000", X"00000000", X"c6589045"),
		(X"4312199a", X"00000000", X"c658dc71"),
		(X"43123333", X"00000000", X"c65928aa"),
		(X"43124ccd", X"00000000", X"c65974f1"),
		(X"43126666", X"00000000", X"c659c145"),
		(X"43128000", X"00000000", X"c65a0da7"),
		(X"4312999a", X"00000000", X"c65a5a16"),
		(X"4312b333", X"00000000", X"c65aa692"),
		(X"4312cccd", X"00000000", X"c65af31c"),
		(X"4312e666", X"00000000", X"c65b3fb3"),
		(X"43130000", X"00000000", X"c65b8c57"),
		(X"4313199a", X"00000000", X"c65bd909"),
		(X"43133333", X"00000000", X"c65c25c8"),
		(X"43134ccd", X"00000000", X"c65c7295"),
		(X"43136666", X"00000000", X"c65cbf6f"),
		(X"43138000", X"00000000", X"c65d0c56"),
		(X"4313999a", X"00000000", X"c65d594b"),
		(X"4313b333", X"00000000", X"c65da64d"),
		(X"4313cccd", X"00000000", X"c65df35c"),
		(X"4313e666", X"00000000", X"c65e4079"),
		(X"43140000", X"00000000", X"45c47ab1"),
		(X"4314199a", X"00000000", X"45c4be49"),
		(X"43143333", X"00000000", X"45c501ed"),
		(X"43144ccd", X"00000000", X"45c5459c"),
		(X"43146666", X"00000000", X"45c58957"),
		(X"43148000", X"00000000", X"45c5cd1e"),
		(X"4314999a", X"00000000", X"45c610f0"),
		(X"4314b333", X"00000000", X"45c654cd"),
		(X"4314cccd", X"00000000", X"45c698b7"),
		(X"4314e666", X"00000000", X"45c6dcac"),
		(X"43150000", X"00000000", X"45c720ac"),
		(X"4315199a", X"00000000", X"45c764b9"),
		(X"43153333", X"00000000", X"45c7a8d0"),
		(X"43154ccd", X"00000000", X"45c7ecf4"),
		(X"43156666", X"00000000", X"45c83123"),
		(X"43158000", X"00000000", X"45c8755e"),
		(X"4315999a", X"00000000", X"45c8b9a4"),
		(X"4315b333", X"00000000", X"45c8fdf6"),
		(X"4315cccd", X"00000000", X"45c94254"),
		(X"4315e666", X"00000000", X"45c986bd"),
		(X"43160000", X"00000000", X"45c9cb32"),
		(X"4316199a", X"00000000", X"45ca0fb2"),
		(X"43163333", X"00000000", X"45ca543e"),
		(X"43164ccd", X"00000000", X"45ca98d6"),
		(X"43166666", X"00000000", X"45cadd79"),
		(X"43168000", X"00000000", X"45cb2228"),
		(X"4316999a", X"00000000", X"45cb66e2"),
		(X"4316b333", X"00000000", X"45cbaba8"),
		(X"4316cccd", X"00000000", X"45cbf07a"),
		(X"4316e666", X"00000000", X"45cc3558"),
		(X"43170000", X"00000000", X"45cc7a40"),
		(X"4317199a", X"00000000", X"45ccbf35"),
		(X"43173333", X"00000000", X"45cd0435"),
		(X"43174ccd", X"00000000", X"45cd4941"),
		(X"43176666", X"00000000", X"45cd8e59"),
		(X"43178000", X"00000000", X"45cdd37c"),
		(X"4317999a", X"00000000", X"45ce18aa"),
		(X"4317b333", X"00000000", X"45ce5de5"),
		(X"4317cccd", X"00000000", X"45cea32b"),
		(X"4317e666", X"00000000", X"45cee87c"),
		(X"43180000", X"00000000", X"46ade78c"),
		(X"4318199a", X"00000000", X"46ae220c"),
		(X"43183333", X"00000000", X"46ae5c95"),
		(X"43184ccd", X"00000000", X"46ae9728"),
		(X"43186666", X"00000000", X"46aed1c5"),
		(X"43188000", X"00000000", X"46af0c6c"),
		(X"4318999a", X"00000000", X"46af471c"),
		(X"4318b333", X"00000000", X"46af81d7"),
		(X"4318cccd", X"00000000", X"46afbc9b"),
		(X"4318e666", X"00000000", X"46aff769"),
		(X"43190000", X"00000000", X"46b03241"),
		(X"4319199a", X"00000000", X"46b06d22"),
		(X"43193333", X"00000000", X"46b0a80e"),
		(X"43194ccd", X"00000000", X"46b0e303"),
		(X"43196666", X"00000000", X"46b11e02"),
		(X"43198000", X"00000000", X"46b1590b"),
		(X"4319999a", X"00000000", X"46b1941e"),
		(X"4319b333", X"00000000", X"46b1cf3b"),
		(X"4319cccd", X"00000000", X"46b20a62"),
		(X"4319e666", X"00000000", X"46b24592"),
		(X"431a0000", X"00000000", X"46b280cc"),
		(X"431a199a", X"00000000", X"46b2bc10"),
		(X"431a3333", X"00000000", X"46b2f75e"),
		(X"431a4ccd", X"00000000", X"46b332b6"),
		(X"431a6666", X"00000000", X"46b36e17"),
		(X"431a8000", X"00000000", X"46b3a982"),
		(X"431a999a", X"00000000", X"46b3e4f8"),
		(X"431ab333", X"00000000", X"46b42077"),
		(X"431acccd", X"00000000", X"46b45bff"),
		(X"431ae666", X"00000000", X"46b49792"),
		(X"431b0000", X"00000000", X"46b4d32f"),
		(X"431b199a", X"00000000", X"46b50ed5"),
		(X"431b3333", X"00000000", X"46b54a85"),
		(X"431b4ccd", X"00000000", X"46b5863f"),
		(X"431b6666", X"00000000", X"46b5c203"),
		(X"431b8000", X"00000000", X"46b5fdd1"),
		(X"431b999a", X"00000000", X"46b639a8"),
		(X"431bb333", X"00000000", X"46b6758a"),
		(X"431bcccd", X"00000000", X"46b6b175"),
		(X"431be666", X"00000000", X"46b6ed6a"),
		(X"431c0000", X"00000000", X"468ff1ee"),
		(X"431c199a", X"00000000", X"46902117"),
		(X"431c3333", X"00000000", X"46905047"),
		(X"431c4ccd", X"00000000", X"46907f7f"),
		(X"431c6666", X"00000000", X"4690aebf"),
		(X"431c8000", X"00000000", X"4690de06"),
		(X"431c999a", X"00000000", X"46910d56"),
		(X"431cb333", X"00000000", X"46913cad"),
		(X"431ccccd", X"00000000", X"46916c0b"),
		(X"431ce666", X"00000000", X"46919b71"),
		(X"431d0000", X"00000000", X"4691cae0"),
		(X"431d199a", X"00000000", X"4691fa55"),
		(X"431d3333", X"00000000", X"469229d3"),
		(X"431d4ccd", X"00000000", X"46925958"),
		(X"431d6666", X"00000000", X"469288e5"),
		(X"431d8000", X"00000000", X"4692b87a"),
		(X"431d999a", X"00000000", X"4692e816"),
		(X"431db333", X"00000000", X"469317ba"),
		(X"431dcccd", X"00000000", X"46934766"),
		(X"431de666", X"00000000", X"4693771a"),
		(X"431e0000", X"00000000", X"4693a6d5"),
		(X"431e199a", X"00000000", X"4693d698"),
		(X"431e3333", X"00000000", X"46940663"),
		(X"431e4ccd", X"00000000", X"46943635"),
		(X"431e6666", X"00000000", X"4694660f"),
		(X"431e8000", X"00000000", X"469495f1"),
		(X"431e999a", X"00000000", X"4694c5db"),
		(X"431eb333", X"00000000", X"4694f5cc"),
		(X"431ecccd", X"00000000", X"469525c5"),
		(X"431ee666", X"00000000", X"469555c6"),
		(X"431f0000", X"00000000", X"469585ce"),
		(X"431f199a", X"00000000", X"4695b5de"),
		(X"431f3333", X"00000000", X"4695e5f6"),
		(X"431f4ccd", X"00000000", X"46961616"),
		(X"431f6666", X"00000000", X"4696463d"),
		(X"431f8000", X"00000000", X"4696766c"),
		(X"431f999a", X"00000000", X"4696a6a3"),
		(X"431fb333", X"00000000", X"4696d6e2"),
		(X"431fcccd", X"00000000", X"46970728"),
		(X"431fe666", X"00000000", X"46973776"),
		(X"43200000", X"00000000", X"c563ccd0"),
		(X"4320199a", X"00000000", X"c5641688"),
		(X"43203333", X"00000000", X"c564604d"),
		(X"43204ccd", X"00000000", X"c564aa1d"),
		(X"43206666", X"00000000", X"c564f3f8"),
		(X"43208000", X"00000000", X"c5653de0"),
		(X"4320999a", X"00000000", X"c56587d4"),
		(X"4320b333", X"00000000", X"c565d1d4"),
		(X"4320cccd", X"00000000", X"c5661bdf"),
		(X"4320e666", X"00000000", X"c56665f7"),
		(X"43210000", X"00000000", X"c566b01a"),
		(X"4321199a", X"00000000", X"c566fa49"),
		(X"43213333", X"00000000", X"c5674485"),
		(X"43214ccd", X"00000000", X"c5678ecc"),
		(X"43216666", X"00000000", X"c567d91f"),
		(X"43218000", X"00000000", X"c568237e"),
		(X"4321999a", X"00000000", X"c5686de9"),
		(X"4321b333", X"00000000", X"c568b860"),
		(X"4321cccd", X"00000000", X"c56902e3"),
		(X"4321e666", X"00000000", X"c5694d71"),
		(X"43220000", X"00000000", X"c569980c"),
		(X"4322199a", X"00000000", X"c569e2b2"),
		(X"43223333", X"00000000", X"c56a2d65"),
		(X"43224ccd", X"00000000", X"c56a7823"),
		(X"43226666", X"00000000", X"c56ac2ed"),
		(X"43228000", X"00000000", X"c56b0dc4"),
		(X"4322999a", X"00000000", X"c56b58a6"),
		(X"4322b333", X"00000000", X"c56ba394"),
		(X"4322cccd", X"00000000", X"c56bee8e"),
		(X"4322e666", X"00000000", X"c56c3994"),
		(X"43230000", X"00000000", X"c56c84a5"),
		(X"4323199a", X"00000000", X"c56ccfc3"),
		(X"43233333", X"00000000", X"c56d1aed"),
		(X"43234ccd", X"00000000", X"c56d6622"),
		(X"43236666", X"00000000", X"c56db164"),
		(X"43238000", X"00000000", X"c56dfcb1"),
		(X"4323999a", X"00000000", X"c56e480b"),
		(X"4323b333", X"00000000", X"c56e9370"),
		(X"4323cccd", X"00000000", X"c56edee1"),
		(X"4323e666", X"00000000", X"c56f2a5e"),
		(X"43240000", X"00000000", X"c6becf85"),
		(X"4324199a", X"00000000", X"c6bf0b35"),
		(X"43243333", X"00000000", X"c6bf46ef"),
		(X"43244ccd", X"00000000", X"c6bf82b2"),
		(X"43246666", X"00000000", X"c6bfbe7e"),
		(X"43248000", X"00000000", X"c6bffa53"),
		(X"4324999a", X"00000000", X"c6c03632"),
		(X"4324b333", X"00000000", X"c6c0721a"),
		(X"4324cccd", X"00000000", X"c6c0ae0c"),
		(X"4324e666", X"00000000", X"c6c0ea07"),
		(X"43250000", X"00000000", X"c6c1260b"),
		(X"4325199a", X"00000000", X"c6c16218"),
		(X"43253333", X"00000000", X"c6c19e2f"),
		(X"43254ccd", X"00000000", X"c6c1da50"),
		(X"43256666", X"00000000", X"c6c21679"),
		(X"43258000", X"00000000", X"c6c252ac"),
		(X"4325999a", X"00000000", X"c6c28ee8"),
		(X"4325b333", X"00000000", X"c6c2cb2e"),
		(X"4325cccd", X"00000000", X"c6c3077c"),
		(X"4325e666", X"00000000", X"c6c343d5"),
		(X"43260000", X"00000000", X"c6c38036"),
		(X"4326199a", X"00000000", X"c6c3bca1"),
		(X"43263333", X"00000000", X"c6c3f915"),
		(X"43264ccd", X"00000000", X"c6c43592"),
		(X"43266666", X"00000000", X"c6c47219"),
		(X"43268000", X"00000000", X"c6c4aea9"),
		(X"4326999a", X"00000000", X"c6c4eb43"),
		(X"4326b333", X"00000000", X"c6c527e6"),
		(X"4326cccd", X"00000000", X"c6c56492"),
		(X"4326e666", X"00000000", X"c6c5a147"),
		(X"43270000", X"00000000", X"c6c5de06"),
		(X"4327199a", X"00000000", X"c6c61ace"),
		(X"43273333", X"00000000", X"c6c657a0"),
		(X"43274ccd", X"00000000", X"c6c6947a"),
		(X"43276666", X"00000000", X"c6c6d15f"),
		(X"43278000", X"00000000", X"c6c70e4c"),
		(X"4327999a", X"00000000", X"c6c74b43"),
		(X"4327b333", X"00000000", X"c6c78843"),
		(X"4327cccd", X"00000000", X"c6c7c54c"),
		(X"4327e666", X"00000000", X"c6c8025f"),
		(X"43280000", X"00000000", X"c6b85be9"),
		(X"4328199a", X"00000000", X"c6b89436"),
		(X"43283333", X"00000000", X"c6b8cc8c"),
		(X"43284ccd", X"00000000", X"c6b904eb"),
		(X"43286666", X"00000000", X"c6b93d52"),
		(X"43288000", X"00000000", X"c6b975c2"),
		(X"4328999a", X"00000000", X"c6b9ae3a"),
		(X"4328b333", X"00000000", X"c6b9e6bb"),
		(X"4328cccd", X"00000000", X"c6ba1f45"),
		(X"4328e666", X"00000000", X"c6ba57d7"),
		(X"43290000", X"00000000", X"c6ba9072"),
		(X"4329199a", X"00000000", X"c6bac915"),
		(X"43293333", X"00000000", X"c6bb01c1"),
		(X"43294ccd", X"00000000", X"c6bb3a75"),
		(X"43296666", X"00000000", X"c6bb7333"),
		(X"43298000", X"00000000", X"c6bbabf8"),
		(X"4329999a", X"00000000", X"c6bbe4c7"),
		(X"4329b333", X"00000000", X"c6bc1d9d"),
		(X"4329cccd", X"00000000", X"c6bc567d"),
		(X"4329e666", X"00000000", X"c6bc8f65"),
		(X"432a0000", X"00000000", X"c6bcc856"),
		(X"432a199a", X"00000000", X"c6bd014f"),
		(X"432a3333", X"00000000", X"c6bd3a51"),
		(X"432a4ccd", X"00000000", X"c6bd735b"),
		(X"432a6666", X"00000000", X"c6bdac6e"),
		(X"432a8000", X"00000000", X"c6bde58a"),
		(X"432a999a", X"00000000", X"c6be1eae"),
		(X"432ab333", X"00000000", X"c6be57db"),
		(X"432acccd", X"00000000", X"c6be9110"),
		(X"432ae666", X"00000000", X"c6beca4e"),
		(X"432b0000", X"00000000", X"c6bf0395"),
		(X"432b199a", X"00000000", X"c6bf3ce4"),
		(X"432b3333", X"00000000", X"c6bf763c"),
		(X"432b4ccd", X"00000000", X"c6bfaf9c"),
		(X"432b6666", X"00000000", X"c6bfe905"),
		(X"432b8000", X"00000000", X"c6c02277"),
		(X"432b999a", X"00000000", X"c6c05bf1"),
		(X"432bb333", X"00000000", X"c6c09573"),
		(X"432bcccd", X"00000000", X"c6c0ceff"),
		(X"432be666", X"00000000", X"c6c10893"),
		(X"432c0000", X"00000000", X"4358ee0b"),
		(X"432c199a", X"00000000", X"435921d4"),
		(X"432c3333", X"00000000", X"435955a3"),
		(X"432c4ccd", X"00000000", X"43598977"),
		(X"432c6666", X"00000000", X"4359bd52"),
		(X"432c8000", X"00000000", X"4359f132"),
		(X"432c999a", X"00000000", X"435a2519"),
		(X"432cb333", X"00000000", X"435a5905"),
		(X"432ccccd", X"00000000", X"435a8cf6"),
		(X"432ce666", X"00000000", X"435ac0ee"),
		(X"432d0000", X"00000000", X"435af4eb"),
		(X"432d199a", X"00000000", X"435b28ee"),
		(X"432d3333", X"00000000", X"435b5cf7"),
		(X"432d4ccd", X"00000000", X"435b9106"),
		(X"432d6666", X"00000000", X"435bc51b"),
		(X"432d8000", X"00000000", X"435bf935"),
		(X"432d999a", X"00000000", X"435c2d55"),
		(X"432db333", X"00000000", X"435c617b"),
		(X"432dcccd", X"00000000", X"435c95a7"),
		(X"432de666", X"00000000", X"435cc9d9"),
		(X"432e0000", X"00000000", X"435cfe10"),
		(X"432e199a", X"00000000", X"435d324d"),
		(X"432e3333", X"00000000", X"435d6690"),
		(X"432e4ccd", X"00000000", X"435d9ad9"),
		(X"432e6666", X"00000000", X"435dcf28"),
		(X"432e8000", X"00000000", X"435e037c"),
		(X"432e999a", X"00000000", X"435e37d6"),
		(X"432eb333", X"00000000", X"435e6c36"),
		(X"432ecccd", X"00000000", X"435ea09c"),
		(X"432ee666", X"00000000", X"435ed508"),
		(X"432f0000", X"00000000", X"435f0979"),
		(X"432f199a", X"00000000", X"435f3df0"),
		(X"432f3333", X"00000000", X"435f726d"),
		(X"432f4ccd", X"00000000", X"435fa6f0"),
		(X"432f6666", X"00000000", X"435fdb78"),
		(X"432f8000", X"00000000", X"43601007"),
		(X"432f999a", X"00000000", X"4360449b"),
		(X"432fb333", X"00000000", X"43607935"),
		(X"432fcccd", X"00000000", X"4360add5"),
		(X"432fe666", X"00000000", X"4360e27a"),
		(X"43300000", X"00000000", X"46cce671"),
		(X"4330199a", X"00000000", X"46cd21f7"),
		(X"43303333", X"00000000", X"46cd5d86"),
		(X"43304ccd", X"00000000", X"46cd991d"),
		(X"43306666", X"00000000", X"46cdd4bd"),
		(X"43308000", X"00000000", X"46ce1066"),
		(X"4330999a", X"00000000", X"46ce4c18"),
		(X"4330b333", X"00000000", X"46ce87d2"),
		(X"4330cccd", X"00000000", X"46cec394"),
		(X"4330e666", X"00000000", X"46ceff60"),
		(X"43310000", X"00000000", X"46cf3b34"),
		(X"4331199a", X"00000000", X"46cf7710"),
		(X"43313333", X"00000000", X"46cfb2f5"),
		(X"43314ccd", X"00000000", X"46cfeee3"),
		(X"43316666", X"00000000", X"46d02ada"),
		(X"43318000", X"00000000", X"46d066d9"),
		(X"4331999a", X"00000000", X"46d0a2e1"),
		(X"4331b333", X"00000000", X"46d0def1"),
		(X"4331cccd", X"00000000", X"46d11b0a"),
		(X"4331e666", X"00000000", X"46d1572c"),
		(X"43320000", X"00000000", X"46d19356"),
		(X"4332199a", X"00000000", X"46d1cf89"),
		(X"43323333", X"00000000", X"46d20bc5"),
		(X"43324ccd", X"00000000", X"46d24809"),
		(X"43326666", X"00000000", X"46d28456"),
		(X"43328000", X"00000000", X"46d2c0ac"),
		(X"4332999a", X"00000000", X"46d2fd0a"),
		(X"4332b333", X"00000000", X"46d33971"),
		(X"4332cccd", X"00000000", X"46d375e1"),
		(X"4332e666", X"00000000", X"46d3b259"),
		(X"43330000", X"00000000", X"46d3eed9"),
		(X"4333199a", X"00000000", X"46d42b63"),
		(X"43333333", X"00000000", X"46d467f5"),
		(X"43334ccd", X"00000000", X"46d4a490"),
		(X"43336666", X"00000000", X"46d4e133"),
		(X"43338000", X"00000000", X"46d51ddf"),
		(X"4333999a", X"00000000", X"46d55a94"),
		(X"4333b333", X"00000000", X"46d59751"),
		(X"4333cccd", X"00000000", X"46d5d417"),
		(X"4333e666", X"00000000", X"46d610e5"),
		(X"43340000", X"00000000", X"46e6668d"),
		(X"4334199a", X"00000000", X"46e6a801"),
		(X"43343333", X"00000000", X"46e6e97f"),
		(X"43344ccd", X"00000000", X"46e72b06"),
		(X"43346666", X"00000000", X"46e76c96"),
		(X"43348000", X"00000000", X"46e7ae30"),
		(X"4334999a", X"00000000", X"46e7efd2"),
		(X"4334b333", X"00000000", X"46e8317e"),
		(X"4334cccd", X"00000000", X"46e87334"),
		(X"4334e666", X"00000000", X"46e8b4f2"),
		(X"43350000", X"00000000", X"46e8f6ba"),
		(X"4335199a", X"00000000", X"46e9388c"),
		(X"43353333", X"00000000", X"46e97a66"),
		(X"43354ccd", X"00000000", X"46e9bc4a"),
		(X"43356666", X"00000000", X"46e9fe37"),
		(X"43358000", X"00000000", X"46ea402d"),
		(X"4335999a", X"00000000", X"46ea822d"),
		(X"4335b333", X"00000000", X"46eac436"),
		(X"4335cccd", X"00000000", X"46eb0648"),
		(X"4335e666", X"00000000", X"46eb4864"),
		(X"43360000", X"00000000", X"46eb8a89"),
		(X"4336199a", X"00000000", X"46ebccb7"),
		(X"43363333", X"00000000", X"46ec0eee"),
		(X"43364ccd", X"00000000", X"46ec512f"),
		(X"43366666", X"00000000", X"46ec9379"),
		(X"43368000", X"00000000", X"46ecd5cc"),
		(X"4336999a", X"00000000", X"46ed1829"),
		(X"4336b333", X"00000000", X"46ed5a8f"),
		(X"4336cccd", X"00000000", X"46ed9cfe"),
		(X"4336e666", X"00000000", X"46eddf77"),
		(X"43370000", X"00000000", X"46ee21f8"),
		(X"4337199a", X"00000000", X"46ee6484"),
		(X"43373333", X"00000000", X"46eea718"),
		(X"43374ccd", X"00000000", X"46eee9b6"),
		(X"43376666", X"00000000", X"46ef2c5d"),
		(X"43378000", X"00000000", X"46ef6f0d"),
		(X"4337999a", X"00000000", X"46efb1c6"),
		(X"4337b333", X"00000000", X"46eff489"),
		(X"4337cccd", X"00000000", X"46f03755"),
		(X"4337e666", X"00000000", X"46f07a2b"),
		(X"43380000", X"00000000", X"45938b01"),
		(X"4338199a", X"00000000", X"4593b3ab"),
		(X"43383333", X"00000000", X"4593dc5b"),
		(X"43384ccd", X"00000000", X"45940511"),
		(X"43386666", X"00000000", X"45942dcd"),
		(X"43388000", X"00000000", X"4594568e"),
		(X"4338999a", X"00000000", X"45947f54"),
		(X"4338b333", X"00000000", X"4594a820"),
		(X"4338cccd", X"00000000", X"4594d0f2"),
		(X"4338e666", X"00000000", X"4594f9c9"),
		(X"43390000", X"00000000", X"459522a6"),
		(X"4339199a", X"00000000", X"45954b89"),
		(X"43393333", X"00000000", X"45957471"),
		(X"43394ccd", X"00000000", X"45959d5f"),
		(X"43396666", X"00000000", X"4595c652"),
		(X"43398000", X"00000000", X"4595ef4b"),
		(X"4339999a", X"00000000", X"4596184a"),
		(X"4339b333", X"00000000", X"4596414e"),
		(X"4339cccd", X"00000000", X"45966a58"),
		(X"4339e666", X"00000000", X"45969368"),
		(X"433a0000", X"00000000", X"4596bc7d"),
		(X"433a199a", X"00000000", X"4596e597"),
		(X"433a3333", X"00000000", X"45970eb7"),
		(X"433a4ccd", X"00000000", X"459737dd"),
		(X"433a6666", X"00000000", X"45976109"),
		(X"433a8000", X"00000000", X"45978a3a"),
		(X"433a999a", X"00000000", X"4597b370"),
		(X"433ab333", X"00000000", X"4597dcac"),
		(X"433acccd", X"00000000", X"459805ee"),
		(X"433ae666", X"00000000", X"45982f36"),
		(X"433b0000", X"00000000", X"45985883"),
		(X"433b199a", X"00000000", X"459881d5"),
		(X"433b3333", X"00000000", X"4598ab2d"),
		(X"433b4ccd", X"00000000", X"4598d48b"),
		(X"433b6666", X"00000000", X"4598fdef"),
		(X"433b8000", X"00000000", X"45992758"),
		(X"433b999a", X"00000000", X"459950c6"),
		(X"433bb333", X"00000000", X"45997a3b"),
		(X"433bcccd", X"00000000", X"4599a3b4"),
		(X"433be666", X"00000000", X"4599cd34"),
		(X"433c0000", X"00000000", X"c6d108d2"),
		(X"433c199a", X"00000000", X"c6d141dd"),
		(X"433c3333", X"00000000", X"c6d17af0"),
		(X"433c4ccd", X"00000000", X"c6d1b40b"),
		(X"433c6666", X"00000000", X"c6d1ed2d"),
		(X"433c8000", X"00000000", X"c6d22657"),
		(X"433c999a", X"00000000", X"c6d25f8a"),
		(X"433cb333", X"00000000", X"c6d298c3"),
		(X"433ccccd", X"00000000", X"c6d2d205"),
		(X"433ce666", X"00000000", X"c6d30b4f"),
		(X"433d0000", X"00000000", X"c6d344a0"),
		(X"433d199a", X"00000000", X"c6d37df9"),
		(X"433d3333", X"00000000", X"c6d3b759"),
		(X"433d4ccd", X"00000000", X"c6d3f0c2"),
		(X"433d6666", X"00000000", X"c6d42a32"),
		(X"433d8000", X"00000000", X"c6d463aa"),
		(X"433d999a", X"00000000", X"c6d49d2a"),
		(X"433db333", X"00000000", X"c6d4d6b2"),
		(X"433dcccd", X"00000000", X"c6d51041"),
		(X"433de666", X"00000000", X"c6d549d9"),
		(X"433e0000", X"00000000", X"c6d58378"),
		(X"433e199a", X"00000000", X"c6d5bd1e"),
		(X"433e3333", X"00000000", X"c6d5f6cd"),
		(X"433e4ccd", X"00000000", X"c6d63083"),
		(X"433e6666", X"00000000", X"c6d66a41"),
		(X"433e8000", X"00000000", X"c6d6a407"),
		(X"433e999a", X"00000000", X"c6d6ddd5"),
		(X"433eb333", X"00000000", X"c6d717aa"),
		(X"433ecccd", X"00000000", X"c6d75188"),
		(X"433ee666", X"00000000", X"c6d78b6d"),
		(X"433f0000", X"00000000", X"c6d7c559"),
		(X"433f199a", X"00000000", X"c6d7ff4e"),
		(X"433f3333", X"00000000", X"c6d8394a"),
		(X"433f4ccd", X"00000000", X"c6d8734f"),
		(X"433f6666", X"00000000", X"c6d8ad5a"),
		(X"433f8000", X"00000000", X"c6d8e76e"),
		(X"433f999a", X"00000000", X"c6d9218a"),
		(X"433fb333", X"00000000", X"c6d95bad"),
		(X"433fcccd", X"00000000", X"c6d995d8"),
		(X"433fe666", X"00000000", X"c6d9d00b"),
		(X"43400000", X"00000000", X"c7098729"),
		(X"4340199a", X"00000000", X"c709abe5"),
		(X"43403333", X"00000000", X"c709d0a5"),
		(X"43404ccd", X"00000000", X"c709f56b"),
		(X"43406666", X"00000000", X"c70a1a35"),
		(X"43408000", X"00000000", X"c70a3f05"),
		(X"4340999a", X"00000000", X"c70a63d9"),
		(X"4340b333", X"00000000", X"c70a88b2"),
		(X"4340cccd", X"00000000", X"c70aad91"),
		(X"4340e666", X"00000000", X"c70ad274"),
		(X"43410000", X"00000000", X"c70af75c"),
		(X"4341199a", X"00000000", X"c70b1c49"),
		(X"43413333", X"00000000", X"c70b413a"),
		(X"43414ccd", X"00000000", X"c70b6631"),
		(X"43416666", X"00000000", X"c70b8b2d"),
		(X"43418000", X"00000000", X"c70bb02d"),
		(X"4341999a", X"00000000", X"c70bd532"),
		(X"4341b333", X"00000000", X"c70bfa3d"),
		(X"4341cccd", X"00000000", X"c70c1f4c"),
		(X"4341e666", X"00000000", X"c70c4460"),
		(X"43420000", X"00000000", X"c70c6979"),
		(X"4342199a", X"00000000", X"c70c8e97"),
		(X"43423333", X"00000000", X"c70cb3ba"),
		(X"43424ccd", X"00000000", X"c70cd8e1"),
		(X"43426666", X"00000000", X"c70cfe0e"),
		(X"43428000", X"00000000", X"c70d233f"),
		(X"4342999a", X"00000000", X"c70d4876"),
		(X"4342b333", X"00000000", X"c70d6db1"),
		(X"4342cccd", X"00000000", X"c70d92f1"),
		(X"4342e666", X"00000000", X"c70db836"),
		(X"43430000", X"00000000", X"c70ddd80"),
		(X"4343199a", X"00000000", X"c70e02cf"),
		(X"43433333", X"00000000", X"c70e2823"),
		(X"43434ccd", X"00000000", X"c70e4d7c"),
		(X"43436666", X"00000000", X"c70e72da"),
		(X"43438000", X"00000000", X"c70e983c"),
		(X"4343999a", X"00000000", X"c70ebda4"),
		(X"4343b333", X"00000000", X"c70ee310"),
		(X"4343cccd", X"00000000", X"c70f0881"),
		(X"4343e666", X"00000000", X"c70f2df7"),
		(X"43440000", X"00000000", X"c623a2b3"),
		(X"4344199a", X"00000000", X"c623cda8"),
		(X"43443333", X"00000000", X"c623f8a2"),
		(X"43444ccd", X"00000000", X"c62423a3"),
		(X"43446666", X"00000000", X"c6244ea8"),
		(X"43448000", X"00000000", X"c62479b4"),
		(X"4344999a", X"00000000", X"c624a4c5"),
		(X"4344b333", X"00000000", X"c624cfdc"),
		(X"4344cccd", X"00000000", X"c624faf8"),
		(X"4344e666", X"00000000", X"c625261a"),
		(X"43450000", X"00000000", X"c6255142"),
		(X"4345199a", X"00000000", X"c6257c6f"),
		(X"43453333", X"00000000", X"c625a7a2"),
		(X"43454ccd", X"00000000", X"c625d2da"),
		(X"43456666", X"00000000", X"c625fe18"),
		(X"43458000", X"00000000", X"c626295c"),
		(X"4345999a", X"00000000", X"c62654a6"),
		(X"4345b333", X"00000000", X"c6267ff5"),
		(X"4345cccd", X"00000000", X"c626ab49"),
		(X"4345e666", X"00000000", X"c626d6a4"),
		(X"43460000", X"00000000", X"c6270204"),
		(X"4346199a", X"00000000", X"c6272d69"),
		(X"43463333", X"00000000", X"c62758d4"),
		(X"43464ccd", X"00000000", X"c6278445"),
		(X"43466666", X"00000000", X"c627afbc"),
		(X"43468000", X"00000000", X"c627db38"),
		(X"4346999a", X"00000000", X"c62806ba"),
		(X"4346b333", X"00000000", X"c6283241"),
		(X"4346cccd", X"00000000", X"c6285dce"),
		(X"4346e666", X"00000000", X"c6288961"),
		(X"43470000", X"00000000", X"c628b4f9"),
		(X"4347199a", X"00000000", X"c628e097"),
		(X"43473333", X"00000000", X"c6290c3b"),
		(X"43474ccd", X"00000000", X"c62937e4"),
		(X"43476666", X"00000000", X"c6296393"),
		(X"43478000", X"00000000", X"c6298f47"),
		(X"4347999a", X"00000000", X"c629bb01"),
		(X"4347b333", X"00000000", X"c629e6c1"),
		(X"4347cccd", X"00000000", X"c62a1287"),
		(X"4347e666", X"00000000", X"c62a3e52"),
		(X"43480000", X"00000000", X"46cf2156"),
		(X"4348199a", X"00000000", X"46cf5646"),
		(X"43483333", X"00000000", X"46cf8b3d"),
		(X"43484ccd", X"00000000", X"46cfc03b"),
		(X"43486666", X"00000000", X"46cff540"),
		(X"43488000", X"00000000", X"46d02a4b"),
		(X"4348999a", X"00000000", X"46d05f5d"),
		(X"4348b333", X"00000000", X"46d09476"),
		(X"4348cccd", X"00000000", X"46d0c996"),
		(X"4348e666", X"00000000", X"46d0febc"),
		(X"43490000", X"00000000", X"46d133e9"),
		(X"4349199a", X"00000000", X"46d1691d"),
		(X"43493333", X"00000000", X"46d19e58"),
		(X"43494ccd", X"00000000", X"46d1d399"),
		(X"43496666", X"00000000", X"46d208e1"),
		(X"43498000", X"00000000", X"46d23e30"),
		(X"4349999a", X"00000000", X"46d27386"),
		(X"4349b333", X"00000000", X"46d2a8e2"),
		(X"4349cccd", X"00000000", X"46d2de46"),
		(X"4349e666", X"00000000", X"46d313af"),
		(X"434a0000", X"00000000", X"46d34920"),
		(X"434a199a", X"00000000", X"46d37e98"),
		(X"434a3333", X"00000000", X"46d3b416"),
		(X"434a4ccd", X"00000000", X"46d3e99b"),
		(X"434a6666", X"00000000", X"46d41f27"),
		(X"434a8000", X"00000000", X"46d454b9"),
		(X"434a999a", X"00000000", X"46d48a53"),
		(X"434ab333", X"00000000", X"46d4bff3"),
		(X"434acccd", X"00000000", X"46d4f59a"),
		(X"434ae666", X"00000000", X"46d52b47"),
		(X"434b0000", X"00000000", X"46d560fc"),
		(X"434b199a", X"00000000", X"46d596b7"),
		(X"434b3333", X"00000000", X"46d5cc79"),
		(X"434b4ccd", X"00000000", X"46d60241"),
		(X"434b6666", X"00000000", X"46d63811"),
		(X"434b8000", X"00000000", X"46d66de7"),
		(X"434b999a", X"00000000", X"46d6a3c4"),
		(X"434bb333", X"00000000", X"46d6d9a7"),
		(X"434bcccd", X"00000000", X"46d70f92"),
		(X"434be666", X"00000000", X"46d74583"),
		(X"434c0000", X"00000000", X"47211fee"),
		(X"434c199a", X"00000000", X"47214855"),
		(X"434c3333", X"00000000", X"472170c0"),
		(X"434c4ccd", X"00000000", X"47219930"),
		(X"434c6666", X"00000000", X"4721c1a5"),
		(X"434c8000", X"00000000", X"4721ea20"),
		(X"434c999a", X"00000000", X"4722129f"),
		(X"434cb333", X"00000000", X"47223b24"),
		(X"434ccccd", X"00000000", X"472263ad"),
		(X"434ce666", X"00000000", X"47228c3c"),
		(X"434d0000", X"00000000", X"4722b4d0"),
		(X"434d199a", X"00000000", X"4722dd69"),
		(X"434d3333", X"00000000", X"47230606"),
		(X"434d4ccd", X"00000000", X"47232ea9"),
		(X"434d6666", X"00000000", X"47235751"),
		(X"434d8000", X"00000000", X"47237ffe"),
		(X"434d999a", X"00000000", X"4723a8b0"),
		(X"434db333", X"00000000", X"4723d167"),
		(X"434dcccd", X"00000000", X"4723fa24"),
		(X"434de666", X"00000000", X"472422e5"),
		(X"434e0000", X"00000000", X"47244bab"),
		(X"434e199a", X"00000000", X"47247477"),
		(X"434e3333", X"00000000", X"47249d47"),
		(X"434e4ccd", X"00000000", X"4724c61d"),
		(X"434e6666", X"00000000", X"4724eef7"),
		(X"434e8000", X"00000000", X"472517d7"),
		(X"434e999a", X"00000000", X"472540bc"),
		(X"434eb333", X"00000000", X"472569a5"),
		(X"434ecccd", X"00000000", X"47259294"),
		(X"434ee666", X"00000000", X"4725bb88"),
		(X"434f0000", X"00000000", X"4725e481"),
		(X"434f199a", X"00000000", X"47260d7f"),
		(X"434f3333", X"00000000", X"47263682"),
		(X"434f4ccd", X"00000000", X"47265f8a"),
		(X"434f6666", X"00000000", X"47268898"),
		(X"434f8000", X"00000000", X"4726b1aa"),
		(X"434f999a", X"00000000", X"4726dac1"),
		(X"434fb333", X"00000000", X"472703de"),
		(X"434fcccd", X"00000000", X"47272cff"),
		(X"434fe666", X"00000000", X"47275625"),
		(X"43500000", X"00000000", X"468abe86"),
		(X"4350199a", X"00000000", X"468ae096"),
		(X"43503333", X"00000000", X"468b02aa"),
		(X"43504ccd", X"00000000", X"468b24c1"),
		(X"43506666", X"00000000", X"468b46dd"),
		(X"43508000", X"00000000", X"468b68fe"),
		(X"4350999a", X"00000000", X"468b8b22"),
		(X"4350b333", X"00000000", X"468bad4b"),
		(X"4350cccd", X"00000000", X"468bcf77"),
		(X"4350e666", X"00000000", X"468bf1a8"),
		(X"43510000", X"00000000", X"468c13dd"),
		(X"4351199a", X"00000000", X"468c3617"),
		(X"43513333", X"00000000", X"468c5854"),
		(X"43514ccd", X"00000000", X"468c7a96"),
		(X"43516666", X"00000000", X"468c9cdc"),
		(X"43518000", X"00000000", X"468cbf26"),
		(X"4351999a", X"00000000", X"468ce174"),
		(X"4351b333", X"00000000", X"468d03c6"),
		(X"4351cccd", X"00000000", X"468d261d"),
		(X"4351e666", X"00000000", X"468d4878"),
		(X"43520000", X"00000000", X"468d6ad6"),
		(X"4352199a", X"00000000", X"468d8d3a"),
		(X"43523333", X"00000000", X"468dafa1"),
		(X"43524ccd", X"00000000", X"468dd20c"),
		(X"43526666", X"00000000", X"468df47c"),
		(X"43528000", X"00000000", X"468e16f0"),
		(X"4352999a", X"00000000", X"468e3968"),
		(X"4352b333", X"00000000", X"468e5be4"),
		(X"4352cccd", X"00000000", X"468e7e64"),
		(X"4352e666", X"00000000", X"468ea0e9"),
		(X"43530000", X"00000000", X"468ec371"),
		(X"4353199a", X"00000000", X"468ee5fe"),
		(X"43533333", X"00000000", X"468f088f"),
		(X"43534ccd", X"00000000", X"468f2b25"),
		(X"43536666", X"00000000", X"468f4dbe"),
		(X"43538000", X"00000000", X"468f705c"),
		(X"4353999a", X"00000000", X"468f92fd"),
		(X"4353b333", X"00000000", X"468fb5a3"),
		(X"4353cccd", X"00000000", X"468fd84d"),
		(X"4353e666", X"00000000", X"468ffafc"),
		(X"43540000", X"00000000", X"c6bf7e4a"),
		(X"4354199a", X"00000000", X"c6bfaca5"),
		(X"43543333", X"00000000", X"c6bfdb07"),
		(X"43544ccd", X"00000000", X"c6c0096e"),
		(X"43546666", X"00000000", X"c6c037da"),
		(X"43548000", X"00000000", X"c6c0664c"),
		(X"4354999a", X"00000000", X"c6c094c4"),
		(X"4354b333", X"00000000", X"c6c0c342"),
		(X"4354cccd", X"00000000", X"c6c0f1c5"),
		(X"4354e666", X"00000000", X"c6c1204d"),
		(X"43550000", X"00000000", X"c6c14edc"),
		(X"4355199a", X"00000000", X"c6c17d6f"),
		(X"43553333", X"00000000", X"c6c1ac09"),
		(X"43554ccd", X"00000000", X"c6c1daa8"),
		(X"43556666", X"00000000", X"c6c2094d"),
		(X"43558000", X"00000000", X"c6c237f7"),
		(X"4355999a", X"00000000", X"c6c266a7"),
		(X"4355b333", X"00000000", X"c6c2955c"),
		(X"4355cccd", X"00000000", X"c6c2c417"),
		(X"4355e666", X"00000000", X"c6c2f2d8"),
		(X"43560000", X"00000000", X"c6c3219e"),
		(X"4356199a", X"00000000", X"c6c3506a"),
		(X"43563333", X"00000000", X"c6c37f3c"),
		(X"43564ccd", X"00000000", X"c6c3ae13"),
		(X"43566666", X"00000000", X"c6c3dcf0"),
		(X"43568000", X"00000000", X"c6c40bd2"),
		(X"4356999a", X"00000000", X"c6c43aba"),
		(X"4356b333", X"00000000", X"c6c469a8"),
		(X"4356cccd", X"00000000", X"c6c4989b"),
		(X"4356e666", X"00000000", X"c6c4c794"),
		(X"43570000", X"00000000", X"c6c4f692"),
		(X"4357199a", X"00000000", X"c6c52596"),
		(X"43573333", X"00000000", X"c6c554a0"),
		(X"43574ccd", X"00000000", X"c6c583af"),
		(X"43576666", X"00000000", X"c6c5b2c4"),
		(X"43578000", X"00000000", X"c6c5e1de"),
		(X"4357999a", X"00000000", X"c6c610fe"),
		(X"4357b333", X"00000000", X"c6c64024"),
		(X"4357cccd", X"00000000", X"c6c66f4f"),
		(X"4357e666", X"00000000", X"c6c69e80"),
		(X"43580000", X"00000000", X"c735d22c"),
		(X"4358199a", X"00000000", X"c735fd55"),
		(X"43583333", X"00000000", X"c7362882"),
		(X"43584ccd", X"00000000", X"c73653b5"),
		(X"43586666", X"00000000", X"c7367eed"),
		(X"43588000", X"00000000", X"c736aa2a"),
		(X"4358999a", X"00000000", X"c736d56c"),
		(X"4358b333", X"00000000", X"c73700b3"),
		(X"4358cccd", X"00000000", X"c7372c00"),
		(X"4358e666", X"00000000", X"c7375751"),
		(X"43590000", X"00000000", X"c73782a8"),
		(X"4359199a", X"00000000", X"c737ae03"),
		(X"43593333", X"00000000", X"c737d964"),
		(X"43594ccd", X"00000000", X"c73804ca"),
		(X"43596666", X"00000000", X"c7383035"),
		(X"43598000", X"00000000", X"c7385ba6"),
		(X"4359999a", X"00000000", X"c738871b"),
		(X"4359b333", X"00000000", X"c738b295"),
		(X"4359cccd", X"00000000", X"c738de15"),
		(X"4359e666", X"00000000", X"c739099a"),
		(X"435a0000", X"00000000", X"c7393523"),
		(X"435a199a", X"00000000", X"c73960b2"),
		(X"435a3333", X"00000000", X"c7398c46"),
		(X"435a4ccd", X"00000000", X"c739b7e0"),
		(X"435a6666", X"00000000", X"c739e37e"),
		(X"435a8000", X"00000000", X"c73a0f21"),
		(X"435a999a", X"00000000", X"c73a3aca"),
		(X"435ab333", X"00000000", X"c73a6677"),
		(X"435acccd", X"00000000", X"c73a922a"),
		(X"435ae666", X"00000000", X"c73abde2"),
		(X"435b0000", X"00000000", X"c73ae99f"),
		(X"435b199a", X"00000000", X"c73b1561"),
		(X"435b3333", X"00000000", X"c73b4128"),
		(X"435b4ccd", X"00000000", X"c73b6cf5"),
		(X"435b6666", X"00000000", X"c73b98c6"),
		(X"435b8000", X"00000000", X"c73bc49d"),
		(X"435b999a", X"00000000", X"c73bf079"),
		(X"435bb333", X"00000000", X"c73c1c59"),
		(X"435bcccd", X"00000000", X"c73c483f"),
		(X"435be666", X"00000000", X"c73c742a"),
		(X"435c0000", X"00000000", X"c6c89e3d"),
		(X"435c199a", X"00000000", X"c6c8cd09"),
		(X"435c3333", X"00000000", X"c6c8fbdc"),
		(X"435c4ccd", X"00000000", X"c6c92ab3"),
		(X"435c6666", X"00000000", X"c6c95990"),
		(X"435c8000", X"00000000", X"c6c98873"),
		(X"435c999a", X"00000000", X"c6c9b75b"),
		(X"435cb333", X"00000000", X"c6c9e649"),
		(X"435ccccd", X"00000000", X"c6ca153c"),
		(X"435ce666", X"00000000", X"c6ca4434"),
		(X"435d0000", X"00000000", X"c6ca7332"),
		(X"435d199a", X"00000000", X"c6caa235"),
		(X"435d3333", X"00000000", X"c6cad13e"),
		(X"435d4ccd", X"00000000", X"c6cb004c"),
		(X"435d6666", X"00000000", X"c6cb2f60"),
		(X"435d8000", X"00000000", X"c6cb5e79"),
		(X"435d999a", X"00000000", X"c6cb8d98"),
		(X"435db333", X"00000000", X"c6cbbcbc"),
		(X"435dcccd", X"00000000", X"c6cbebe6"),
		(X"435de666", X"00000000", X"c6cc1b15"),
		(X"435e0000", X"00000000", X"c6cc4a49"),
		(X"435e199a", X"00000000", X"c6cc7983"),
		(X"435e3333", X"00000000", X"c6cca8c2"),
		(X"435e4ccd", X"00000000", X"c6ccd807"),
		(X"435e6666", X"00000000", X"c6cd0751"),
		(X"435e8000", X"00000000", X"c6cd36a1"),
		(X"435e999a", X"00000000", X"c6cd65f6"),
		(X"435eb333", X"00000000", X"c6cd9551"),
		(X"435ecccd", X"00000000", X"c6cdc4b1"),
		(X"435ee666", X"00000000", X"c6cdf417"),
		(X"435f0000", X"00000000", X"c6ce2382"),
		(X"435f199a", X"00000000", X"c6ce52f2"),
		(X"435f3333", X"00000000", X"c6ce8268"),
		(X"435f4ccd", X"00000000", X"c6ceb1e3"),
		(X"435f6666", X"00000000", X"c6cee164"),
		(X"435f8000", X"00000000", X"c6cf10eb"),
		(X"435f999a", X"00000000", X"c6cf4076"),
		(X"435fb333", X"00000000", X"c6cf7008"),
		(X"435fcccd", X"00000000", X"c6cf9f9e"),
		(X"435fe666", X"00000000", X"c6cfcf3a"),
		(X"43600000", X"00000000", X"46a72736"),
		(X"4360199a", X"00000000", X"46a74d54"),
		(X"43603333", X"00000000", X"46a77375"),
		(X"43604ccd", X"00000000", X"46a7999b"),
		(X"43606666", X"00000000", X"46a7bfc6"),
		(X"43608000", X"00000000", X"46a7e5f5"),
		(X"4360999a", X"00000000", X"46a80c28"),
		(X"4360b333", X"00000000", X"46a8325f"),
		(X"4360cccd", X"00000000", X"46a8589b"),
		(X"4360e666", X"00000000", X"46a87edb"),
		(X"43610000", X"00000000", X"46a8a520"),
		(X"4361199a", X"00000000", X"46a8cb69"),
		(X"43613333", X"00000000", X"46a8f1b6"),
		(X"43614ccd", X"00000000", X"46a91807"),
		(X"43616666", X"00000000", X"46a93e5d"),
		(X"43618000", X"00000000", X"46a964b8"),
		(X"4361999a", X"00000000", X"46a98b16"),
		(X"4361b333", X"00000000", X"46a9b179"),
		(X"4361cccd", X"00000000", X"46a9d7e0"),
		(X"4361e666", X"00000000", X"46a9fe4c"),
		(X"43620000", X"00000000", X"46aa24bc"),
		(X"4362199a", X"00000000", X"46aa4b30"),
		(X"43623333", X"00000000", X"46aa71a9"),
		(X"43624ccd", X"00000000", X"46aa9826"),
		(X"43626666", X"00000000", X"46aabea7"),
		(X"43628000", X"00000000", X"46aae52d"),
		(X"4362999a", X"00000000", X"46ab0bb7"),
		(X"4362b333", X"00000000", X"46ab3245"),
		(X"4362cccd", X"00000000", X"46ab58d8"),
		(X"4362e666", X"00000000", X"46ab7f6f"),
		(X"43630000", X"00000000", X"46aba60a"),
		(X"4363199a", X"00000000", X"46abccaa"),
		(X"43633333", X"00000000", X"46abf34e"),
		(X"43634ccd", X"00000000", X"46ac19f6"),
		(X"43636666", X"00000000", X"46ac40a3"),
		(X"43638000", X"00000000", X"46ac6754"),
		(X"4363999a", X"00000000", X"46ac8e0a"),
		(X"4363b333", X"00000000", X"46acb4c4"),
		(X"4363cccd", X"00000000", X"46acdb82"),
		(X"4363e666", X"00000000", X"46ad0244"),
		(X"43640000", X"00000000", X"4749b8b0"),
		(X"4364199a", X"00000000", X"4749e5f2"),
		(X"43643333", X"00000000", X"474a1339"),
		(X"43644ccd", X"00000000", X"474a4086"),
		(X"43646666", X"00000000", X"474a6dd7"),
		(X"43648000", X"00000000", X"474a9b2e"),
		(X"4364999a", X"00000000", X"474ac889"),
		(X"4364b333", X"00000000", X"474af5ea"),
		(X"4364cccd", X"00000000", X"474b2350"),
		(X"4364e666", X"00000000", X"474b50bb"),
		(X"43650000", X"00000000", X"474b7e2b"),
		(X"4365199a", X"00000000", X"474baba0"),
		(X"43653333", X"00000000", X"474bd91a"),
		(X"43654ccd", X"00000000", X"474c0699"),
		(X"43656666", X"00000000", X"474c341d"),
		(X"43658000", X"00000000", X"474c61a6"),
		(X"4365999a", X"00000000", X"474c8f35"),
		(X"4365b333", X"00000000", X"474cbcc8"),
		(X"4365cccd", X"00000000", X"474cea61"),
		(X"4365e666", X"00000000", X"474d17fe"),
		(X"43660000", X"00000000", X"474d45a1"),
		(X"4366199a", X"00000000", X"474d7349"),
		(X"43663333", X"00000000", X"474da0f6"),
		(X"43664ccd", X"00000000", X"474dcea7"),
		(X"43666666", X"00000000", X"474dfc5e"),
		(X"43668000", X"00000000", X"474e2a1a"),
		(X"4366999a", X"00000000", X"474e57dc"),
		(X"4366b333", X"00000000", X"474e85a2"),
		(X"4366cccd", X"00000000", X"474eb36d"),
		(X"4366e666", X"00000000", X"474ee13d"),
		(X"43670000", X"00000000", X"474f0f13"),
		(X"4367199a", X"00000000", X"474f3ced"),
		(X"43673333", X"00000000", X"474f6acd"),
		(X"43674ccd", X"00000000", X"474f98b1"),
		(X"43676666", X"00000000", X"474fc69b"),
		(X"43678000", X"00000000", X"474ff48a"),
		(X"4367999a", X"00000000", X"4750227e"),
		(X"4367b333", X"00000000", X"47505077"),
		(X"4367cccd", X"00000000", X"47507e75"),
		(X"4367e666", X"00000000", X"4750ac78"),
		(X"43680000", X"00000000", X"470877c9"),
		(X"4368199a", X"00000000", X"470895dc"),
		(X"43683333", X"00000000", X"4708b3f2"),
		(X"43684ccd", X"00000000", X"4708d20c"),
		(X"43686666", X"00000000", X"4708f028"),
		(X"43688000", X"00000000", X"47090e48"),
		(X"4368999a", X"00000000", X"47092c6c"),
		(X"4368b333", X"00000000", X"47094a92"),
		(X"4368cccd", X"00000000", X"470968bc"),
		(X"4368e666", X"00000000", X"470986ea"),
		(X"43690000", X"00000000", X"4709a51a"),
		(X"4369199a", X"00000000", X"4709c34e"),
		(X"43693333", X"00000000", X"4709e186"),
		(X"43694ccd", X"00000000", X"4709ffc0"),
		(X"43696666", X"00000000", X"470a1dfe"),
		(X"43698000", X"00000000", X"470a3c3f"),
		(X"4369999a", X"00000000", X"470a5a84"),
		(X"4369b333", X"00000000", X"470a78cc"),
		(X"4369cccd", X"00000000", X"470a9717"),
		(X"4369e666", X"00000000", X"470ab565"),
		(X"436a0000", X"00000000", X"470ad3b7"),
		(X"436a199a", X"00000000", X"470af20c"),
		(X"436a3333", X"00000000", X"470b1064"),
		(X"436a4ccd", X"00000000", X"470b2ec0"),
		(X"436a6666", X"00000000", X"470b4d1f"),
		(X"436a8000", X"00000000", X"470b6b81"),
		(X"436a999a", X"00000000", X"470b89e7"),
		(X"436ab333", X"00000000", X"470ba850"),
		(X"436acccd", X"00000000", X"470bc6bc"),
		(X"436ae666", X"00000000", X"470be52c"),
		(X"436b0000", X"00000000", X"470c039f"),
		(X"436b199a", X"00000000", X"470c2215"),
		(X"436b3333", X"00000000", X"470c408e"),
		(X"436b4ccd", X"00000000", X"470c5f0b"),
		(X"436b6666", X"00000000", X"470c7d8b"),
		(X"436b8000", X"00000000", X"470c9c0f"),
		(X"436b999a", X"00000000", X"470cba95"),
		(X"436bb333", X"00000000", X"470cd91f"),
		(X"436bcccd", X"00000000", X"470cf7ad"),
		(X"436be666", X"00000000", X"470d163e"),
		(X"436c0000", X"00000000", X"c67c63da"),
		(X"436c199a", X"00000000", X"c67c9ad2"),
		(X"436c3333", X"00000000", X"c67cd1d0"),
		(X"436c4ccd", X"00000000", X"c67d08d3"),
		(X"436c6666", X"00000000", X"c67d3fdd"),
		(X"436c8000", X"00000000", X"c67d76ec"),
		(X"436c999a", X"00000000", X"c67dae02"),
		(X"436cb333", X"00000000", X"c67de51e"),
		(X"436ccccd", X"00000000", X"c67e1c3f"),
		(X"436ce666", X"00000000", X"c67e5367"),
		(X"436d0000", X"00000000", X"c67e8a94"),
		(X"436d199a", X"00000000", X"c67ec1c8"),
		(X"436d3333", X"00000000", X"c67ef901"),
		(X"436d4ccd", X"00000000", X"c67f3041"),
		(X"436d6666", X"00000000", X"c67f6786"),
		(X"436d8000", X"00000000", X"c67f9ed2"),
		(X"436d999a", X"00000000", X"c67fd623"),
		(X"436db333", X"00000000", X"c68006bd"),
		(X"436dcccd", X"00000000", X"c680226c"),
		(X"436de666", X"00000000", X"c6803e1e"),
		(X"436e0000", X"00000000", X"c68059d2"),
		(X"436e199a", X"00000000", X"c680758a"),
		(X"436e3333", X"00000000", X"c6809145"),
		(X"436e4ccd", X"00000000", X"c680ad02"),
		(X"436e6666", X"00000000", X"c680c8c3"),
		(X"436e8000", X"00000000", X"c680e487"),
		(X"436e999a", X"00000000", X"c681004d"),
		(X"436eb333", X"00000000", X"c6811c17"),
		(X"436ecccd", X"00000000", X"c68137e3"),
		(X"436ee666", X"00000000", X"c68153b3"),
		(X"436f0000", X"00000000", X"c6816f86"),
		(X"436f199a", X"00000000", X"c6818b5b"),
		(X"436f3333", X"00000000", X"c681a734"),
		(X"436f4ccd", X"00000000", X"c681c30f"),
		(X"436f6666", X"00000000", X"c681deee"),
		(X"436f8000", X"00000000", X"c681facf"),
		(X"436f999a", X"00000000", X"c68216b4"),
		(X"436fb333", X"00000000", X"c682329b"),
		(X"436fcccd", X"00000000", X"c6824e86"),
		(X"436fe666", X"00000000", X"c6826a74"),
		(X"43700000", X"00000000", X"c7581e19"),
		(X"4370199a", X"00000000", X"c7584c43"),
		(X"43703333", X"00000000", X"c7587a72"),
		(X"43704ccd", X"00000000", X"c758a8a6"),
		(X"43706666", X"00000000", X"c758d6df"),
		(X"43708000", X"00000000", X"c759051d"),
		(X"4370999a", X"00000000", X"c7593360"),
		(X"4370b333", X"00000000", X"c75961a8"),
		(X"4370cccd", X"00000000", X"c7598ff4"),
		(X"4370e666", X"00000000", X"c759be46"),
		(X"43710000", X"00000000", X"c759ec9c"),
		(X"4371199a", X"00000000", X"c75a1af8"),
		(X"43713333", X"00000000", X"c75a4958"),
		(X"43714ccd", X"00000000", X"c75a77be"),
		(X"43716666", X"00000000", X"c75aa628"),
		(X"43718000", X"00000000", X"c75ad497"),
		(X"4371999a", X"00000000", X"c75b030b"),
		(X"4371b333", X"00000000", X"c75b3184"),
		(X"4371cccd", X"00000000", X"c75b6002"),
		(X"4371e666", X"00000000", X"c75b8e85"),
		(X"43720000", X"00000000", X"c75bbd0d"),
		(X"4372199a", X"00000000", X"c75beb9a"),
		(X"43723333", X"00000000", X"c75c1a2b"),
		(X"43724ccd", X"00000000", X"c75c48c2"),
		(X"43726666", X"00000000", X"c75c775d"),
		(X"43728000", X"00000000", X"c75ca5fe"),
		(X"4372999a", X"00000000", X"c75cd4a3"),
		(X"4372b333", X"00000000", X"c75d034d"),
		(X"4372cccd", X"00000000", X"c75d31fd"),
		(X"4372e666", X"00000000", X"c75d60b1"),
		(X"43730000", X"00000000", X"c75d8f6a"),
		(X"4373199a", X"00000000", X"c75dbe28"),
		(X"43733333", X"00000000", X"c75deceb"),
		(X"43734ccd", X"00000000", X"c75e1bb3"),
		(X"43736666", X"00000000", X"c75e4a80"),
		(X"43738000", X"00000000", X"c75e7951"),
		(X"4373999a", X"00000000", X"c75ea828"),
		(X"4373b333", X"00000000", X"c75ed704"),
		(X"4373cccd", X"00000000", X"c75f05e4"),
		(X"4373e666", X"00000000", X"c75f34ca"),
		(X"43740000", X"00000000", X"c72d7e5a"),
		(X"4374199a", X"00000000", X"c72da2d1"),
		(X"43743333", X"00000000", X"c72dc74b"),
		(X"43744ccd", X"00000000", X"c72debc9"),
		(X"43746666", X"00000000", X"c72e104b"),
		(X"43748000", X"00000000", X"c72e34d1"),
		(X"4374999a", X"00000000", X"c72e595b"),
		(X"4374b333", X"00000000", X"c72e7de8"),
		(X"4374cccd", X"00000000", X"c72ea279"),
		(X"4374e666", X"00000000", X"c72ec70e"),
		(X"43750000", X"00000000", X"c72eeba7"),
		(X"4375199a", X"00000000", X"c72f1044"),
		(X"43753333", X"00000000", X"c72f34e5"),
		(X"43754ccd", X"00000000", X"c72f5989"),
		(X"43756666", X"00000000", X"c72f7e31"),
		(X"43758000", X"00000000", X"c72fa2dd"),
		(X"4375999a", X"00000000", X"c72fc78d"),
		(X"4375b333", X"00000000", X"c72fec41"),
		(X"4375cccd", X"00000000", X"c73010f8"),
		(X"4375e666", X"00000000", X"c73035b4"),
		(X"43760000", X"00000000", X"c7305a73"),
		(X"4376199a", X"00000000", X"c7307f36"),
		(X"43763333", X"00000000", X"c730a3fd"),
		(X"43764ccd", X"00000000", X"c730c8c8"),
		(X"43766666", X"00000000", X"c730ed96"),
		(X"43768000", X"00000000", X"c7311269"),
		(X"4376999a", X"00000000", X"c731373f"),
		(X"4376b333", X"00000000", X"c7315c19"),
		(X"4376cccd", X"00000000", X"c73180f7"),
		(X"4376e666", X"00000000", X"c731a5d8"),
		(X"43770000", X"00000000", X"c731cabe"),
		(X"4377199a", X"00000000", X"c731efa7"),
		(X"43773333", X"00000000", X"c7321494"),
		(X"43774ccd", X"00000000", X"c7323985"),
		(X"43776666", X"00000000", X"c7325e7a"),
		(X"43778000", X"00000000", X"c7328373"),
		(X"4377999a", X"00000000", X"c732a86f"),
		(X"4377b333", X"00000000", X"c732cd70"),
		(X"4377cccd", X"00000000", X"c732f274"),
		(X"4377e666", X"00000000", X"c733177c"),
		(X"43780000", X"00000000", X"46162c53"),
		(X"4378199a", X"00000000", X"46164b22"),
		(X"43783333", X"00000000", X"461669f5"),
		(X"43784ccd", X"00000000", X"461688ca"),
		(X"43786666", X"00000000", X"4616a7a3"),
		(X"43788000", X"00000000", X"4616c67f"),
		(X"4378999a", X"00000000", X"4616e55e"),
		(X"4378b333", X"00000000", X"46170440"),
		(X"4378cccd", X"00000000", X"46172326"),
		(X"4378e666", X"00000000", X"4617420e"),
		(X"43790000", X"00000000", X"461760fa"),
		(X"4379199a", X"00000000", X"46177fe9"),
		(X"43793333", X"00000000", X"46179edb"),
		(X"43794ccd", X"00000000", X"4617bdd0"),
		(X"43796666", X"00000000", X"4617dcc8"),
		(X"43798000", X"00000000", X"4617fbc4"),
		(X"4379999a", X"00000000", X"46181ac3"),
		(X"4379b333", X"00000000", X"461839c4"),
		(X"4379cccd", X"00000000", X"461858c9"),
		(X"4379e666", X"00000000", X"461877d1"),
		(X"437a0000", X"00000000", X"461896dd"),
		(X"437a199a", X"00000000", X"4618b5eb"),
		(X"437a3333", X"00000000", X"4618d4fd"),
		(X"437a4ccd", X"00000000", X"4618f412"),
		(X"437a6666", X"00000000", X"4619132a"),
		(X"437a8000", X"00000000", X"46193245"),
		(X"437a999a", X"00000000", X"46195163"),
		(X"437ab333", X"00000000", X"46197084"),
		(X"437acccd", X"00000000", X"46198fa9"),
		(X"437ae666", X"00000000", X"4619aed1"),
		(X"437b0000", X"00000000", X"4619cdfb"),
		(X"437b199a", X"00000000", X"4619ed2a"),
		(X"437b3333", X"00000000", X"461a0c5b"),
		(X"437b4ccd", X"00000000", X"461a2b8f"),
		(X"437b6666", X"00000000", X"461a4ac7"),
		(X"437b8000", X"00000000", X"461a6a01"),
		(X"437b999a", X"00000000", X"461a893f"),
		(X"437bb333", X"00000000", X"461aa880"),
		(X"437bcccd", X"00000000", X"461ac7c4"),
		(X"437be666", X"00000000", X"461ae70c"),
		(X"437c0000", X"00000000", X"476367cc"),
		(X"437c199a", X"00000000", X"476395f6"),
		(X"437c3333", X"00000000", X"4763c424"),
		(X"437c4ccd", X"00000000", X"4763f257"),
		(X"437c6666", X"00000000", X"4764208f"),
		(X"437c8000", X"00000000", X"47644ecb"),
		(X"437c999a", X"00000000", X"47647d0c"),
		(X"437cb333", X"00000000", X"4764ab51"),
		(X"437ccccd", X"00000000", X"4764d99c"),
		(X"437ce666", X"00000000", X"476507eb"),
		(X"437d0000", X"00000000", X"4765363e"),
		(X"437d199a", X"00000000", X"47656497"),
		(X"437d3333", X"00000000", X"476592f4"),
		(X"437d4ccd", X"00000000", X"4765c155"),
		(X"437d6666", X"00000000", X"4765efbc"),
		(X"437d8000", X"00000000", X"47661e27"),
		(X"437d999a", X"00000000", X"47664c97"),
		(X"437db333", X"00000000", X"47667b0b"),
		(X"437dcccd", X"00000000", X"4766a984"),
		(X"437de666", X"00000000", X"4766d802"),
		(X"437e0000", X"00000000", X"47670685"),
		(X"437e199a", X"00000000", X"4767350c"),
		(X"437e3333", X"00000000", X"47676398"),
		(X"437e4ccd", X"00000000", X"47679228"),
		(X"437e6666", X"00000000", X"4767c0bd"),
		(X"437e8000", X"00000000", X"4767ef57"),
		(X"437e999a", X"00000000", X"47681df6"),
		(X"437eb333", X"00000000", X"47684c99"),
		(X"437ecccd", X"00000000", X"47687b41"),
		(X"437ee666", X"00000000", X"4768a9ee"),
		(X"437f0000", X"00000000", X"4768d89f"),
		(X"437f199a", X"00000000", X"47690755"),
		(X"437f3333", X"00000000", X"47693610"),
		(X"437f4ccd", X"00000000", X"476964cf"),
		(X"437f6666", X"00000000", X"47699393"),
		(X"437f8000", X"00000000", X"4769c25c"),
		(X"437f999a", X"00000000", X"4769f12a"),
		(X"437fb333", X"00000000", X"476a1ffc"),
		(X"437fcccd", X"00000000", X"476a4ed2"),
		(X"437fe666", X"00000000", X"476a7dae"),
		(X"00000000", X"00000000", X"00000000"),
		(X"40a00000", X"00000000", X"41caf2cf"),
		(X"41200000", X"41caf2cf", X"42372cc1"),
		(X"41700000", X"42372cc1", X"c2e609da"),
		(X"41a00000", X"c2e609da", X"c35ddff1"),
		(X"41c80000", X"c35ddff1", X"4342f327"),
		(X"41f00000", X"4342f327", X"4489c109"),
		(X"420c0000", X"4489c109", X"44cce4da"),
		(X"42200000", X"44cce4da", X"426cdb73"),
		(X"42340000", X"426cdb73", X"c4806e00"),
		(X"42480000", X"c4806e00", X"418e2444"),
		(X"425c0000", X"418e2444", X"453dc196"),
		(X"42700000", X"453dc196", X"4501b82e"),
		(X"42820000", X"4501b82e", X"c4f24334"),
		(X"428c0000", X"c4f24334", X"c5afcc91"),
		(X"42960000", X"c5afcc91", X"c5969764"),
		(X"42a00000", X"c5969764", X"441b6f71"),
		(X"42aa0000", X"441b6f71", X"442e0de2"),
		(X"42b40000", X"442e0de2", X"c5bd3a19"),
		(X"42be0000", X"c5bd3a19", X"c65e5ada"),
		(X"42c80000", X"c65e5ada", X"c5cf8d86"),
		(X"42d20000", X"c5cf8d86", X"4579cafe"),
		(X"42dc0000", X"4579cafe", X"45e9dfff"),
		(X"42e60000", X"45e9dfff", X"c489de00"),
		(X"42f00000", X"c489de00", X"c5dbdb9e"),
		(X"42fa0000", X"c5dbdb9e", X"44b7a8b0"),
		(X"43020000", X"44b7a8b0", X"4690048b"),
		(X"43070000", X"4690048b", X"46dd7990"),
		(X"430c0000", X"46dd7990", X"460cdbb6"),
		(X"43110000", X"460cdbb6", X"c5917b6f"),
		(X"43160000", X"c5917b6f", X"44e13f0c"),
		(X"431b0000", X"44e13f0c", X"46c2e71f"),
		(X"43200000", X"46c2e71f", X"46a66d85"),
		(X"43250000", X"46a66d85", X"c555c42d"),
		(X"432a0000", X"c555c42d", X"c6d780db"),
		(X"432f0000", X"c6d780db", X"c6d5c2c8"),
		(X"43340000", X"c6d5c2c8", X"45051e27"),
		(X"43390000", X"45051e27", X"45d7b1ba"),
		(X"433e0000", X"45d7b1ba", X"c69f9709"),
		(X"43430000", X"c69f9709", X"c75da905"),
		(X"43480000", X"c75da905", X"c6ec30b4"),
		(X"434d0000", X"c6ec30b4", X"463271d7"),
		(X"43520000", X"463271d7", X"46e6a3c2"),
		(X"43570000", X"46e6a3c2", X"4586b4c1"),
		(X"435c0000", X"4586b4c1", X"c6a6f10c"),
		(X"43610000", X"c6a6f10c", X"435a09d0"),
		(X"43660000", X"435a09d0", X"474e1fab"),
		(X"436b0000", X"474e1fab", X"47ad11a5"),
		(X"43700000", X"47ad11a5", X"47020530"),
		(X"43750000", X"47020530", X"c63399dc"),
		(X"437a0000", X"c63399dc", X"c4d817f7"),
		(X"437f0000", X"c4d817f7", X"476217df")
	);
END PACKAGE fp_mult_data_pak;
