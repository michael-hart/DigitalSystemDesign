LIBRARY IEEE;
LIBRARY IEEE_proposed;

USE IEEE.std_logic_1164.ALL;
USE IEEE_proposed.fixed_pkg.ALL;

PACKAGE cos_data_pak IS

	-- Define data types array
	TYPE data_t_rec IS
		RECORD
      		data, result : sfixed(1 DOWNTO -22);
		END RECORD;
	TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;
	
	-- Define actual data
	CONSTANT data : data_t := (
		(X"000000", X"400000"),
		(X"0066F1", X"3FFFAD"),
		(X"00CDE3", X"3FFEB4"),
		(X"0134D4", X"3FFD16"),
		(X"019BC6", X"3FFAD3"),
		(X"0202B7", X"3FF7EA"),
		(X"0269A9", X"3FF45B"),
		(X"02D09B", X"3FF027"),
		(X"03378C", X"3FEB4E"),
		(X"039E7E", X"3FE5CF"),
		(X"04056F", X"3FDFAB"),
		(X"046C61", X"3FD8E2"),
		(X"04D353", X"3FD173"),
		(X"053A44", X"3FC95F"),
		(X"05A136", X"3FC0A7"),
		(X"060827", X"3FB749"),
		(X"066F19", X"3FAD47"),
		(X"06D60B", X"3FA29F"),
		(X"073CFC", X"3F9753"),
		(X"07A3EE", X"3F8B63"),
		(X"080ADF", X"3F7ECE"),
		(X"0871D1", X"3F7195"),
		(X"08D8C2", X"3F63B8"),
		(X"093FB4", X"3F5537"),
		(X"09A6A6", X"3F4611"),
		(X"0A0D97", X"3F3649"),
		(X"0A7489", X"3F25DC"),
		(X"0ADB7A", X"3F14CD"),
		(X"0B426C", X"3F031A"),
		(X"0BA95E", X"3EF0C4"),
		(X"0C104F", X"3EDDCB"),
		(X"0C7741", X"3ECA2F"),
		(X"0CDE32", X"3EB5F1"),
		(X"0D4524", X"3EA111"),
		(X"0DAC16", X"3E8B8F"),
		(X"0E1307", X"3E756B"),
		(X"0E79F9", X"3E5EA5"),
		(X"0EE0EA", X"3E473E"),
		(X"0F47DC", X"3E2F36"),
		(X"0FAECD", X"3E168D"),
		(X"1015BF", X"3DFD44"),
		(X"107CB1", X"3DE35A"),
		(X"10E3A2", X"3DC8D0"),
		(X"114A94", X"3DADA6"),
		(X"11B185", X"3D91DC"),
		(X"121877", X"3D7573"),
		(X"127F69", X"3D586B"),
		(X"12E65A", X"3D3AC5"),
		(X"134D4C", X"3D1C80"),
		(X"13B43D", X"3CFD9D"),
		(X"141B2F", X"3CDE1C"),
		(X"148221", X"3CBDFD"),
		(X"14E912", X"3C9D42"),
		(X"155004", X"3C7BE9"),
		(X"15B6F5", X"3C59F4"),
		(X"161DE7", X"3C3763"),
		(X"1684D8", X"3C1437"),
		(X"16EBCA", X"3BF06E"),
		(X"1752BC", X"3BCC0B"),
		(X"17B9AD", X"3BA70D"),
		(X"18209F", X"3B8175"),
		(X"188790", X"3B5B42"),
		(X"18EE82", X"3B3477"),
		(X"195574", X"3B0D11"),
		(X"19BC65", X"3AE514"),
		(X"1A2357", X"3ABC7D"),
		(X"1A8A48", X"3A934F"),
		(X"1AF13A", X"3A6989"),
		(X"1B582C", X"3A3F2D"),
		(X"1BBF1D", X"3A1439"),
		(X"1C260F", X"39E8AF"),
		(X"1C8D00", X"39BC90"),
		(X"1CF3F2", X"398FDB"),
		(X"1D5AE4", X"396291"),
		(X"1DC1D5", X"3934B2"),
		(X"1E28C7", X"390640"),
		(X"1E8FB8", X"38D73A"),
		(X"1EF6AA", X"38A7A1"),
		(X"1F5D9B", X"387775"),
		(X"1FC48D", X"3846B7"),
		(X"202B7F", X"381568"),
		(X"209270", X"37E388"),
		(X"20F962", X"37B117"),
		(X"216053", X"377E16"),
		(X"21C745", X"374A85"),
		(X"222E37", X"371665"),
		(X"229528", X"36E1B7"),
		(X"22FC1A", X"36AC7B"),
		(X"23630B", X"3676B1"),
		(X"23C9FD", X"36405A"),
		(X"2430EF", X"360977"),
		(X"2497E0", X"35D209"),
		(X"24FED2", X"359A0F"),
		(X"2565C3", X"35618A"),
		(X"25CCB5", X"35287B"),
		(X"2633A6", X"34EEE3"),
		(X"269A98", X"34B4C2"),
		(X"27018A", X"347A18"),
		(X"27687B", X"343EE6"),
		(X"27CF6D", X"34032E"),
		(X"28365E", X"33C6EF"),
		(X"289D50", X"338A2A"),
		(X"290442", X"334CDF"),
		(X"296B33", X"330F10"),
		(X"29D225", X"32D0BD"),
		(X"2A3916", X"3291E6"),
		(X"2AA008", X"32528C"),
		(X"2B06FA", X"3212B0"),
		(X"2B6DEB", X"31D253"),
		(X"2BD4DD", X"319175"),
		(X"2C3BCE", X"315016"),
		(X"2CA2C0", X"310E38"),
		(X"2D09B1", X"30CBDB"),
		(X"2D70A3", X"308900"),
		(X"2DD795", X"3045A7"),
		(X"2E3E86", X"3001D1"),
		(X"2EA578", X"2FBD7F"),
		(X"2F0C69", X"2F78B2"),
		(X"2F735B", X"2F336A"),
		(X"2FDA4D", X"2EEDA7"),
		(X"30413E", X"2EA76C"),
		(X"30A830", X"2E60B7"),
		(X"310F21", X"2E198B"),
		(X"317613", X"2DD1E7"),
		(X"31DD05", X"2D89CC"),
		(X"3243F6", X"2D413C"),
		(X"32AAE8", X"2CF837"),
		(X"3311D9", X"2CAEBE"),
		(X"3378CB", X"2C64D0"),
		(X"33DFBD", X"2C1A70"),
		(X"3446AE", X"2BCF9E"),
		(X"34ADA0", X"2B845B"),
		(X"351491", X"2B38A7"),
		(X"357B83", X"2AEC83"),
		(X"35E274", X"2A9FF0"),
		(X"364966", X"2A52EF"),
		(X"36B058", X"2A0580"),
		(X"371749", X"29B7A4"),
		(X"377E3B", X"29695D"),
		(X"37E52C", X"291AAA"),
		(X"384C1E", X"28CB8D"),
		(X"38B310", X"287C07"),
		(X"391A01", X"282C18"),
		(X"3980F3", X"27DBC1"),
		(X"39E7E4", X"278B03"),
		(X"3A4ED6", X"2739DE"),
		(X"3AB5C8", X"26E854"),
		(X"3B1CB9", X"269665"),
		(X"3B83AB", X"264413"),
		(X"3BEA9C", X"25F15D"),
		(X"3C518E", X"259E46"),
		(X"3CB87F", X"254ACD"),
		(X"3D1F71", X"24F6F3"),
		(X"3D8663", X"24A2BA"),
		(X"3DED54", X"244E22"),
		(X"3E5446", X"23F92C"),
		(X"3EBB37", X"23A3D9"),
		(X"3F2229", X"234E2A"),
		(X"3F891B", X"22F81F"),
		(X"3FF00C", X"22A1BB"),
		(X"4056FE", X"224AFC"),
		(X"40BDEF", X"21F3E5"),
		(X"4124E1", X"219C76"),
		(X"418BD3", X"2144AF"),
		(X"41F2C4", X"20EC93"),
		(X"4259B6", X"209422"),
		(X"42C0A7", X"203B5C"),
		(X"432799", X"1FE243"),
		(X"438E8A", X"1F88D8"),
		(X"43F57C", X"1F2F1B"),
		(X"445C6E", X"1ED50D"),
		(X"44C35F", X"1E7AAF"),
		(X"452A51", X"1E2003"),
		(X"459142", X"1DC509"),
		(X"45F834", X"1D69C1"),
		(X"465F26", X"1D0E2E"),
		(X"46C617", X"1CB24F"),
		(X"472D09", X"1C5626"),
		(X"4793FA", X"1BF9B4"),
		(X"47FAEC", X"1B9CF9"),
		(X"4861DE", X"1B3FF7"),
		(X"48C8CF", X"1AE2AF"),
		(X"492FC1", X"1A8521"),
		(X"4996B2", X"1A274E"),
		(X"49FDA4", X"19C938"),
		(X"4A6496", X"196ADE"),
		(X"4ACB87", X"190C44"),
		(X"4B3279", X"18AD68"),
		(X"4B996A", X"184E4C"),
		(X"4C005C", X"17EEF2"),
		(X"4C674D", X"178F5A"),
		(X"4CCE3F", X"172F85"),
		(X"4D3531", X"16CF73"),
		(X"4D9C22", X"166F27"),
		(X"4E0314", X"160EA1"),
		(X"4E6A05", X"15ADE1"),
		(X"4ED0F7", X"154CEA"),
		(X"4F37E9", X"14EBBB"),
		(X"4F9EDA", X"148A57"),
		(X"5005CC", X"1428BD"),
		(X"506CBD", X"13C6EF"),
		(X"50D3AF", X"1364EE"),
		(X"513AA1", X"1302BA"),
		(X"51A192", X"12A056"),
		(X"520884", X"123DC1"),
		(X"526F75", X"11DAFD"),
		(X"52D667", X"11780B"),
		(X"533D58", X"1114EC"),
		(X"53A44A", X"10B1A0"),
		(X"540B3C", X"104E29"),
		(X"54722D", X"0FEA88"),
		(X"54D91F", X"0F86BE"),
		(X"554010", X"0F22CC"),
		(X"55A702", X"0EBEB3"),
		(X"560DF4", X"0E5A73"),
		(X"5674E5", X"0DF60F"),
		(X"56DBD7", X"0D9186"),
		(X"5742C8", X"0D2CDA"),
		(X"57A9BA", X"0CC80C"),
		(X"5810AC", X"0C631D"),
		(X"58779D", X"0BFE0E"),
		(X"58DE8F", X"0B98E0"),
		(X"594580", X"0B3393"),
		(X"59AC72", X"0ACE2A"),
		(X"5A1363", X"0A68A5"),
		(X"5A7A55", X"0A0305"),
		(X"5AE147", X"099D4B"),
		(X"5B4838", X"093779"),
		(X"5BAF2A", X"08D18E"),
		(X"5C161B", X"086B8C"),
		(X"5C7D0D", X"080575"),
		(X"5CE3FF", X"079F49"),
		(X"5D4AF0", X"073909"),
		(X"5DB1E2", X"06D2B7"),
		(X"5E18D3", X"066C53"),
		(X"5E7FC5", X"0605DE"),
		(X"5EE6B7", X"059F5A"),
		(X"5F4DA8", X"0538C7"),
		(X"5FB49A", X"04D227"),
		(X"601B8B", X"046B7A"),
		(X"60827D", X"0404C2"),
		(X"60E96F", X"039DFF"),
		(X"615060", X"033733"),
		(X"61B752", X"02D05F"),
		(X"621E43", X"026984"),
		(X"628535", X"0202A2"),
		(X"62EC26", X"019BBB"),
		(X"635318", X"0134D0"),
		(X"63BA0A", X"00CDE1"),
		(X"6420FB", X"0066F1")
	);
END PACKAGE cos_data_pak;
