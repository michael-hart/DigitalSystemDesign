��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F��J>�����>�����HU�k;�� �[�+?�w)݁)��>7Ý�4�B#�"u�%��R9�*2�	φ�v&�f�UxJ�%�����OOL�mF4O0��%�O6?][��W5Ff�i�]�E҅u#��Vg�n�����g9�#���>rh�W&��zCu�M��{����,l6�`I��3����
X�	�@�#��꘲t�}p�ũ�g���.�pæ�dbB�:�`�(8����Q���E�m5���[\[��Z�Xe���z��e�ّ̀�4��'͐??�r���4U��e|{��s�_
���^��5���ЉS�u^R��r	
 K�Ԓ#tO���?�M�ΟuD�(}�G���|E�,n���;��"�z���+�rW�t�ǟ��[�z���Q��Ƈ�b]e}s�;�H�:��(�=����ݺ�����)%����j�⽾I���G6
�<=h��/�[m�S�\I�.4�A�1��S�S��h$��Mj�1�~�P|ul�P�,hM����R2��U�&tˀ.?���9i|������u��F_8�����-�'zx8�~�$	�	+��D\ߍ�b�+/n�f i��O>U�9���mx�������V�K�`?2_�ĥ�3?@A�ʺ*��P �j�C�
����ï��b�A����[���GE��\
���k:
�@�fv6�xR��G��� +�U�.?�T�:y4�_,��7�&��!J�+9?[X��b�1�#���l��;�l���@�7��-�c�)��(�E��V|��i�P/��0��9���E��bQgb
�fYR�E���Do5�����6�r��"�Ҝ��9�=�N���5�Wؒ4��P�bЊ&x�`
'�97^�(9�!W���Dxp@p-/��0Iﴓ8�Y���v-qk��;�Ң7ժ��ٲ?������TH�A���o~��pI��<C�@}|ل1�ў%hz�&��-p�n5�,I�)3�����*�}{�.�O� qI�naG���"0Bσƥ�pl?[� ���,.χcFP��&�?uP��
����������K�,��hXJ��Q��^�M����ϕ��j��#�2��~e�.�Al�Y�1�dY����&p@��>�� 0Θ�2�<�j��S��Z�6G_fo�]7���j�RQ:D���(�՝j���Yo�*�0��cr�}��B��H|ƃ�K1��c-�V�$u�Ɗª��Lo��v0�ƍ���M�m藗���V#����*�Jx�zYr?M�H�>SLL�Xx�$��80�Bd�W�kX}�n��L4�qq��{`�_+\��Yd��}Gi��X}=�Z�tj��^��0	Zu_}�;E*� �{�g�kMK�Z��-T�&���"��OKi�Q(�������ŨrΧw���|l굩mw�޳2�( R�}ׄ�([��Ao�:��VY\\4��fȑ���cSJ�Y�f���-V�3�<�;��hxf�����Z���}���3W�{_�c�)b�S�_m)#���{�c�hb^��)�����`�VG��X՝�>)f)�K����n�I�f��Of���">ږl�{�Deb,��(d?}y���S)j@���$ �7��R_��,�b
5�+�5O��9�c����+������?�+�A�1���vxPƜ��ay�d	�1 1������Ry:����EıD�uz�~���~<WӃz�l��K���h��r�-�z'�?�$aF�?��"ޝ���X���� �R [��z8գN Z�s�D�u	����P���ʜ+~"���H>�u�3A+�1�# ��|�J�ݔ,
M2+��\YC�O5��d��u�{"���,?ؤ��w�7*��;D���"��>wi����D�]�r��,�1B~Ĉ�� �#�y��\����
��Q���4[�J����G��\����_~e��  m��o�/;��;���`u�����w����K��6U���pL`�w{���ޕU6Ɖ�Jv�x����� ~��d�����C� ���>�Y��l�Sx���p5mUT����E=��n�@�)���`J���23����(y�݃���)vW	���YQʰ�Ģ�Ci�Zb�I��|�m�!Y�({� �$�MF"�(NÞ��F��?n�s�QG�І��9��:�����v��� ��ۺv;Y5¼��ྜྷ��}I�H8Z���*q�'{d\ ��.HA���k.��eRA���}��ل�w�^^_~�vk�V(�����#�xcz�R[������@��Z��Nߕi�DDv��k�Ӑ���s�v�2�ְ�(|�CS���T\Ç��h_?憸��J�-�z��0H�ʰlv��-�4��,����(M���:v�_5�y��*�MTIx��EPIη��3�1.���;��z�a�Ʀ5�AaDk�Q�?�B%��\Ζ��ę�
n�ǧ�����3E��c�Qzz��%��E���M-i��L�ka|��C�'�n��@��N�M��[)�2ЖMx�C��̰��=�ߚ$��XЦ9�yסD~"+�3���McK�.a��4%�77f\�����A��WQK3��;8#�WX�T;3y�y� ��|�o�����+��rV����M��'��U��f�cd�uH�}� ��2�c�g�-�Hm{Pܓ��h=�$/���Jy&s�����]e��s�G�k��sk/�R��VKk����X}��뒽!�����U�x["��
9+̗"8ޙ���;V�:�4���P�SU�Lk�ϖR�P ����@�/�K�.f�t�vJ|Q͡/U�j��V�O���s�I\-��=˸g
ۼ3�k����]��F<e�e<uO���A��6��	9��ݵ;��|6����w�������i@l�pP�� ֎����[$E��7$RJ���3�T���x�Gl�Gx~e�w[s*5��3��0B�/fL��eDd'�8Kg� ������*p��0?���95F�j��3���G��p���;�,��D���z���)�i��]��ڇ=�Y_������S5.a� ę��%�ٷ�,��D���!����5֩	�^��Y�ć� E�cI����e�MS[-�ZEK��NDk-�g�t�ؖ��১�����1��-����?�#$����	?A���0pN�u���QD����.����Cn�xm���>����/�0��_d��%�s�>�[��Lj��'8�ʎ:���ӵ�QEg����籟.�A4H��ThY�V�5��N����L��0�ۺA�
�d"L���T�+�#���D�βGM�V�i�h�a�@���Z<��d/�|�]�&��9��
J�u�����>kh��}
�iTڗM!߽�@z����J�ؖ:��Z0ƃ�H�G�.�pV�j*��K��@�Z��U�T��CO�_a� �����}~?ԏ\Mj��Ƥ��k����D��t2�/hݭ+��kHat�5X�����E��t��d�|�)Q���E�\��p��<�BV�����%�֩����E�}bS�y_z/S5c�.s�h?�.�dU���}�!�,N]O����6{y��� �r1 ��/���֖q���<��M$Dk����ϖN�ɮ��+�?�C�-���:�뽉��R��`�`-S�"j�4����Q���R�_���X��I��)�-�2U|�ʼ�����q`.T����W�s���Oz�}�?G5�@��".�PxB�=R$�$����_��(6��]�zuZ���2~�p���|� ׂ�0��<�`��#��EWi�_~�����0�RY�y���
��jGw����D�]L�xH�W��ڟ�Az�9e$8�,U�� ����R��<�B4��t���ԲJ���hqk�s`"v���"o&3<�,~Y��D
c��Dw�xB#�ZaP�C�Y�����[��Ӄ���M�#�a_���W0W���#��1E�#��]���q���D2T�ք"������� �xP&�C�0_gq�/(����7~>3��Ex�Z5��	?�?#���LA�b���{�ڋ�C���O�R\{
�!H01��_�q�qsP����t�!�:$ ir�ķ��R�?�=��+��`�fP�,����l"j��EYm>3Vu���g��پ �ҍ&��S0wM]X���۝�(/�.t��9�f�=�R��ӂC'�ڷSH��5�X��La)��C�!G��N[���j�⇌�3v�ϫ��(�� ��"�����<{%y�y��3�в�kq��t�ª�
s4�e엧虏�c���j�_�!a����ʛm#0|��3��G� ]U?`����O��GI�">F�1̚��N�d�F��xUt�}����`���9���'z���,t�>��,B�{��ULǞT���q����Ѩ��x��ܓ�:.P��1DXӫ���j1���I7^.��28s92N�lHH}e���D|��lJ�c�ސ�yJX����µ�y��r���6;��F����~ f}��Z����c,�5�9D�.�-��1���*��651)�;��H�Ȃ>��t�3��M�����Vs5t��[�wr|���+���H��˄��f��.���N�Tin���*����?(�sC�������v^o���p,)q/^�?��ޒU�D�n���v�5)�!�&e>��rrOb���,rz�j���QO�%��)#j�n�I����jځ��2�����`�~Ȟ?��e��(�!������@m�.����U�\��� O�j֨�c�yȡ	Eg��C�ļ�q��x��c ��)D����>�}#���z��6�������6O?��T�7�5�S�|��+[��`��!�~��[��J9Lg�d�9 ��׍;�	u�ᴮka��|M��9���d=D�?R�2��@թFcL}�\���8XOAl+��)K"�TF���UWs���S6N���M1UG|1�x���-��7:_)hsv�D��G�SCȈf׮����u�8�=�H- ��E�L�9K�I�
��p�����5���j]�5$C'�oQ�}�qN�����PY�tL���%�_8K��ڨq�T�ץ�-�;�,u����I���5
�6B�������lO�i��'�\c���TC��l7�Iy���U�鼸�!H4�m�zX���'�a���(\���Y#�:��9�M/��R�8y�o��jSS�lW;��*ݺur�cFȁ��zؔF) Hߥ-)�.���5�gQ��xq��Y�Yޗ��_�;}��zQ��-&.��M����*�[���r��M �)��RLЕ�~���U���R�!.��b�۸a�=h��n%i��N��T����Aѳ�c�v9���l�'g�7�`M/�D�����2/hH�k��f����Jp<U�W�����b�_N�^'*�?�G/�!n�������؊�g����_��O�RK��,G�O1!�b��,hreG���2 q���[����(��f��1�3{�i���t��{����=_	&/��5Aό$��óS.�8��r*��Y���K}��^���"�H��Yr��i�j4-��Sc�d���L�����@��RB�����%��kef)z��qJ���w�X�#`����Z'�a��Y��Ղ��>�+Y=��I����czx�=�2�6�;
������)IH.r\�J��˯۽]8V��j8K3�dS�*<2�@d$G5��i����v���2cQuY�i�g ZC���T%�d�����*�	8���Y�|L)q0ByЀA�M�~�u��Bр�F��;;��Yf����h�13,������D�'
&�"L����ጃ�
"��ף_Ob4�Єi~�b>Q<�.���F��v�>�>��t�,ĺr?�-�Z>�.e��V�AM[A���<�Q��qZ�������@J94��j��>Q������&<�m�n����Λ���?6X��3���
ǻIxB��Rf��X�"�y���,๛�>7p[d�9�{В�4���W�d�[��فKh�hĢ�.e�9"[`E��9�̪�H�/�e���]О�aW;�������.�Xc�a��@��2��o	u�B�"���"7��]��d�?�J�Vu,TI<'��F_ZU:H/(<��*���u�'d|�y&qJJ��/]�E��v�c�x�u��-C����&?m�u~h�Es�f����+������pK���^��nS�û�(��	h����`�x�*h*W��&�0��
K�z��?\�^�� �Ï�ϕsD��ٛ��!Y�l��[_�@7�_�Èo����t*��3[�]�ė\{2+q#QY���3HX&���o��-�qW
8�h��c9�ҵ;�^��C`�T~��h5�/��<�e�K���כ7O]�CzM}DU>6D�±���J���'�����>��r_\��_�� �Vr�&i�۹���n�'�S��NC`��q$���ǌg2![��	`���������IqWj��eu���T~Ĕ/�A�PP_�*�[��p��WG�4"#YL�ɜ��é����G��<����	��S�Y�T�.q���̓p��Uǎɟ���������p��C�͇��Ρ�	�ꩯ��o%D�s�t$@�tK�G7����x>��m�qʮ\�i۳<�.س�+'>�|EOU�_��3���mw6`��4ñ�}�yǶ��m,;��d�ֵ:���9���Փ��B,s�uIYfP����|�����i��t�5��k�9��%�^�A���E��i���3��5�b�C7�����v�˽�V�O;�hHa�A�ܥ�[�TZ
X�v��]��ݺ���P��ZcB�0�D��<�o�/_���t�T��*�X�:X���B0b����;���x8�eK�>��5�/�Rys�
�ű�&�P�P�I'9R�Ye�d���v��p7�
?t��W٦�g�%̓�wR� 3�)/�+�揋7�@� �b��s�wa��A�M�⤕,+]�y�V�'��BqF�ȿ\1��(@�wI��׼O�w_@T&��������0��(��-�Պ�ҡ�밁��`�!V��=�k\����y�~8�7s�&l\�xϡY>c��'�l�;
���LQ��	�bz���R>\c�Kr5DJ���P8�/�ΐ[��z8%'��O'ZZ�"X��7��
�;��54`�(��b�`7��-����,��+�Q-��#�<l���%Y|��3BH�ǿ&D&�񔿳o��(7R�/���&�]Ж��cz����ULtu�<��E���?�}�ت����BJ�9tŇP�[�Xh!��M۹�쯅p��������"ӟx��l��;%^',�m�÷\�i^3�
*����5�`G��t�>�������=f�j6��7��"��xv5r��&�,�.�̷B��?i��b���0���9o�����F:g����V�w��+�YMGhۣQ����'4��_2�����;{�F�~(e*{�A�lc'|����
T�� T�|��{�HxT�bm42���(����O�IL�W圎��_�t4�B�P9�/�O�9�'�ǁY9�j{�7����v�e{��3X�y���<d�(]i��@L���e�ɼ��@�k�*�f�y�$�����a���f�� �8���1�aF�!@�E!w⾶}��:?�U����|8���"��D�1 ��<���E�F�>��<�d�����	�Z��7�w`6*5�]K�����#� ^���[e3��ϟ���1�M�c9ܕ�_왐 ����g+��ב�ml�:PE�ʯޚ��=�A����.��.���w�,:�kZ�N$W��
�0Lώ����g���T���)+u�����Au{m�w�o�c���5�ƖG{-��r8��lk���rz�C�����:�\R�$
~�Jp��AFH�3���ͥ@����a��c¶+ "������:�|u�_ZpN���Y���&Q�6_����ZH�z��'�L��	k[����U	  w�^��G����E�r#���#pm_ͮ3*�BM�8f���$ohǩ�b��-4���u�����7:����QGZ��5�]�c����Q��ޝV��Y$�/�-dR��7åA��}����L������ ��U��Ɍ�ܮ#��-&�W	;
�DS����`�sL��oi�:�|��!Ǚ+(
��g
ͥ��7N�Q��Nhz�|{��+r(ԃ����+�9��l�H�a�!
Y��7��}�&�;�{�N%/��*�=��Nn߲���tD}I;�2K@�NWm'F�6`6��|3Bn�!Hd���?���Q�� ��&I��C�Rx���P:�N�L��k��Oo%��U4W�w)�:}i�O�G��g9��qd鎣0�N3��p ��o�������	{bBr;�Ҧ�.�U'd��Sp�(h* ����E)p!t�S��D!���6��O�6��))��q����hJX�#�~�	��AY��a8>J��?�S�a�?�"	ӡ��ێL�x�~�9.���tR��K�� N�`�ۭ!�]_����������Ƴ$ʗ�-��Hϥ���`?�R58��tE_<m��7	��W��5�^���ܛC�UA�kx�y*���"(V�> �0o��	�{�̕�)R :4�^.݄�T��.xs�*	:�3�_��]�bޏ����/"ܰz� ��؂�=�,x��:�
�-�&�i����M;����;�0�����n�w��<[�Jl/#�u���u��
�U%d�����C�L�6މ������zJ wR1m侪�c+x'�z}m�!
.&���r�b��jbQD��K���S`��إ�dh��>��4+e�0���UZdz-�'3y���* �Mb��Fb�飳��9�q�@�Ň�:�7��nD���3W�C2++}j�J�;:{&���?���3hY�\��%�Cd̓��]�l��JPd[Y�0r�ǵ�����}�:��(ї�A&�6�m0�i�Ѻ�lqvZ���^`A����<<JM>�.�ό��
nl|�7(���@w���O�w��b5D������q����L��� *�v��aK �l��ݥ�	��n+��)d}Qǲ�P��,��Rd��� �Y$(
�^�wcqðS!Z����𳉍��[+������7��Cm����KR�������t���v�5۩9Q�g���(�����"�X(�or�9�M��/����(j��y��D"ȫi��O��u����
�����)~]ia��	�t�f}�ذ�Ĵ��-��6^ZoGNO�8ვ�����I��Mԏ�(Nˬ��E�a�>�y܆-?�0��{��b�r�=seIv�#"�\x����Zˊ;x<n例l���9�D�al\����k�^�%�5�����Qw֎���7\�"/[���e� ����q�9F��:�%��9��1 *�I��uXAh�ʭM�ѵ�ன���eZ���n�|[��"�Gs@���]����>�6<�����O��a,�_����n=�-������>ڕ�7�p���ɯ@�vX�.B{"�c'��G���8��������  �e����S)�9�2η8�i�T�-d%��|	���;]�SaV�%B�Ӆ*-/���L0���m�h2�K�
� �Ї_=C���ǫ��3%h���gт~P�5�q��\��[��N���2_'�E��۔�8"@��SK�Q}Νo�t�q!����Lk���!
nO̘���qv{�� �~Fʧ�p��xIX$�7�v��j:\,N�2
�?�]�T�~�������Z%��:Tǅ��>+	wq�������&I�����4	�o���m�|��T��w�"�f�"z%T�ێ�����֬&!8y'�����=�2(����j@0|���=������j>�tl׻`з<�{Ɛ`�c��s���Vm�tZh�ش7"�T���K������,9�k���?�Z:卭�Κ�m�?���~����.��u�K�3�~��(K�����Y"L���)���d���G��y�C�'C�}9���oz�ɭ�(N5�j��o��e��ׂ�_����Xg�#>U[7�\�>��� ������pQ@�V�o�9��J�sK#�NPh[R����:s5�	�iB!c��M��D�o>�vΩs�t<�]<E/JčL���2� �3;M@E���(�
c���\�:bW:����v���*u=7���3�v�Dx�J��_��'Y̌��t�Kz�5�J?������I*�I�%ݚJ�qB���ZW�\����W����J�pl�����p�\q�1�&�o�D���>"�yr�o�G�ǥ�,x������G�t��qVi|��'u�&� ��ABF�<�%af&y��^��,��yn��0-?�����~���e����?��*DN�;.{�n�.A.x�T��Z��>���t��Y�Xo�߻�]F!�`�z`ͥYߌ, �:��{;�P2(����-�`�1lC�.��7p�(�Hx�'��x�L>���*)Os5̷��䳨n�vٔ(�]��#�el�R�i�¶����u�%o*��A_�&��H8&�/V���X_k�2?�V���+3���m��-�����u�ز��ZW4�p�Am�V�=�~��/F����
�,̟iE��e�cM�%�v�,U9������ZN+�e+��  r���>)��X���Vm|!`)P@�Zobڤ@��ۛ6�%9p���D����%?��F��/����7*q�xʦKTU��U�8�hk�a�#Ï�O�,�-��FX�ځ��f�[k�-7�xS�-���~�9[Ɵ{X`�el_����_�wȯ "5�^�ߩ+d�*�����Ō��!�P�����ԣ�Ŝ���Bb���I6��C�Z�J����k�Y���L�e���������t����\e�E�H>`N��[�)�t�͎t���R���K�X�-/6G��p%�=� �Z׆!�aܵ���5Ns����s�徸̃
*y����Bw�`�����.��MEI>f��T~:uH��	q8~��ӗC[�'�1�|���l�
�h��uV�;��xǊ>�qa�b�x��r��y�:�%��ڄ�͋�^�=���
w7�>�w��0�J��<��S\'Hkr��C|��,+q� x���<U��n5b4dtl���yO���a��8px�"�q�s1X�yV�0�E�N@ˉ`��4���mi9љ�P���ɨ	�3��|�<�|��uyV>�LHHk�|B�$C��Y6>]��?�x����5?Y�y,�џ�Y�؄�
U���߫���%-����KgȞ�A�ub�P�˶R*�?���P:=��9Q�$U��(��}��2�#!QRaNKNڮ��I�Т)��j+�6��α�;�T�M�Z��;�I�����}0�R�O>d�E0ں8�^���/��48`^6.FjC��N��{M�P��>>q�zӁ�'�J��������i>)��0�d�ME$)w����R����1Vot?���5}r�l�^��8d��JYw	Cǂ���c�ן�K�5lr�����j�}�.K(����'��~�ę�����t���?�z0�A����W�G��y�� ㌳ ~���b�
�u��*����U����������[�E�������50S��~���3���4�N����O��I>S�3iZU	7�̦4ՠT�E��}
s_2��X;�fn�y�!3��{y�,,�����@��l��{U)����3X�n侭�u�Ss;+8�!�}����)�u��`�R��Q	�����:l&�́k��+�1�V�c�@n��H��ݾ�&�l�-(Gwy�<����C��vj��b0�Z��)��x�Q�"��W���T���0�p�������}�=���yXÐ������^�+���8>@���I���C��S=|Km�e#V]o����b��O�~W�=�ه��}RJ4���%oY�d��oב%H���q=�� ���B�C�)���i��zu2�ߨ�眒�-a�-�B5-�ѼN��c-���W'��-R��z}s��3muC��ǘ�[��{��VOB8���Ȼ��B�$�:�΀��/�`��!AtS$�|yl�}A�h�-۱�H&<��*�(*2^�\Y$���`�����+�j0f���1D:���9\�����w��Z�'.ej��ؓ�~^�M�D1�9^��=�vI��K��֏��A�R2Hw�&�Q�f@�`0$ ]z�B^��������{��JD�׍r��n͓Y˿�I�ֵZ7k*4�߱�a�OUL�J�]�)��ݪ ֍�xL�	�z�FHn�V�ýe�;y�X�򝡹����SE�����B�����#q�Ah`��m�[`;�~���MX��:�Ԕ'Ha��:y�����=�h'�ɘ��T���@�p���7i�S�L��x��4���@����8�k��FU � ���,��:o{8{�ll.뫥�?�]�y}{��!�xYa�,sNi
���1���p�'�A�wz����u�����ǖ�.���s��%8�l���ua��Ȣ��sK�I���Q �ʽ�j���Ey+�p^�ruyuC�7��f�m*ޞ+b%�%���߫>��FM�ߨS��8�PA\�K�9�8w��e'���@^��1*������N��7Maz�+��z�B6��9p΁��
1E��`��&_wy���K�>�}ƚ��ؤI����ivk�t�T��l�����a�!�B���q�\v���/��ވ�1\��%l�gq��������l*H/�&${w=S���W���Ĩ˝z�, �(A��*=��~��d�-�����X�Ϻ��`�`C	���7$[� Ɠ��D��Ƅ�S}e(?��ae۲
��x+����4'T�_N�����ܨ|�,�#��M��_*��6�}�9�]�w��4�A ��q>���w����3�u�&T���)i������T�0c�W�m���D���RT��x�zY�a4K�SXW�Ρ��G�k� �UiE�	p3�N�q�Lgq=���
f|O��m�7��E�g��f�bIL��xj=4uƟ��$L8)8����㸓����F	`>eo���f�ǳFH���7�|�C����y�駎ң�����o�v���������U��;�nKgF����)1�5c�룆�{��	�t-�F����֘u��2'ω���{~NԨ�"^��nh6-��3ñ
����U$!l[��E8$f�x�C�@��.�j}k؉��X঑�T� �}�M�뤀��1b����T?�oQr���W/�*�;1���u����#���K2�3D�ӷR�=�(���9�>QԘ�vK�/5;�`(z� 	X4{9!��>�W=ɻ�u��S]�wR���w�90���.:,B'��n�F��[ņ���-��T����$�Wm%`�#�W����"*flv�a��90��T�>C\�t�:��R}�ܞ4ʉ�cmT��4O�Dw�dhТi���x����<��N2�@/�:��X@�QZ�g�����á�J�䶅�]�B��:�YU��3����%U%={������1~d`C�ş?Z�5UȊs*xD�L����0�c� �O��_az�Jxd�=jQ�q�ؗ���ꃓ5⡢|�A4�2��3$IBȘ�w����U�K��$������1�F������t�������(֝ ��?L�{�l:^��7�iO��2'�X;0���$L�4��Q�SqB��|��Ƌn_4�oXx�C�K��C	�M�rE�Cs��eQ|E"��3�8��B P�3HE� ��
�8Z0���7u#A?[�^:a}��1�h�O��4�]0���F�]-X���h!z͐:�%�o,֣W�O�3j�&p"�H�y]o����Ɇ���,%���= �|޴I�M��b���T���8�c�u�`��`Rj�?=�|�"L�Y@Zy�=��,�=lt�d,#\�UhF�Cz��\+�r��EV{���P��Ʌ=��5)5�8C!�����o{���O�i l�-�J��7�:�(%T�Y�zl��8o[���<Ȯd�A3�m6�]���3�ط��܄�yA8A��)5�?�zH�
$�>{�����i/eHTS����j��]����k�-Oz� �U��A׆X��>�y3�����z>�0�UR�y�R�C_Ջ�0�AE�Q�A&�O�3hd�:����|��zr\w���!V�X�sXY�%���
�����f띛ᓶ� �E�ֆ��ǩ櫙��z�?�	f)ò<����8��y�dRٞ[�f;߀*�<���oe֤gq��SиIlC�Z��&�ď}	�`�h$�Y�G
>��uL}i�b��ˎ�4���	>OR����S�Gh�u>�?I=�XP�ʮ�D���3�b�����S�.p4�!1�]�'��Nj!�zǮ`�"��;�������u��ir)�m�P(�kt-ԅw�2g�k���t�?Ӆ�Ap�;���pZ�Z
VA��H[0�3w�i?��6{ݤ�5��w����D��7�8��w������B\X2�Oq�5(n~�4֛�Ҏ~vw��9�P�jx\مm���w%�ڙ���������6���F_p��������R$�>��k�ܱ�DD1� C�IU#ے����Q���b�0�z��p�ˬ��"����qn�Y�;D#�Y,/¼f���� ��ʒ�!Ovd�U�C�1��w�yw�'8#5m��G�m�a�D֟�e���6c7p�l���vUt8MG ��̠hk��V��ӌ��6-+״>Y���dI���whv7<҈�bf�M�*5��saa*;FS�pGٞ�rL��䐢q�s9  ��ەGt�,�26|� ��n�?���F���K�X?-|��|nM]��\�ؑ��y�m��娞�pd~?!;5�1�$h5~a��*�+}&���F=cK��I��K�;��(J)�e�۰V��AF��:�F{z�R[Z��#?Ļ�A"���F(�A�bu��T��M"�^�{��\J ����tI%���:�(D�'�/��@V���$�Ys�|)\�;g�P�S�4@�� ���%�["j{��>��mw_g
��\�#Y#e�%ڬ����}�σė���>������m�
����}+��2
0pFM�फ़��<y�73c�B����&zk����
�)� ⪉=�}�/܃� �FskSchɬi��0�:9uD�'S8� ��>�>�o{�q_Z���Lg��<�j:?i-T�f4�k�%�TLR�!�[v.x]u��4����ǈ�b)��<t�9=�_9�hB�����7�R���THm�Mf~�LQ���E��i��t���a[����R��m*]�2�Q��PO D��z����16�p��<��YŭkSF$��o��R�����ȶ+'�Sҩ"�K���\�	�'(���{��)��;�Ɇ��ұe(F�z�"(��N!�kS)�sXa�!���OXt��ԡ����y�����8�}�0�����0�nJ'>>�6J�ڂ�_�� �V�b�Rjhv�O+�0cu�Z�;���`�6&֟�H���Z}?�,�D�/��Ó`S� L�D��u6��B
-�,�@j��,a��i�j��L�c��;t}o�Ts��!Q*͌c����!7� �^�i�9�A��bַ�N�r�;�)��P���%�X�C���z(�*re�i����W_?��G�*�^�v�������؍c,�Nu
<�E�LbF�eo�2o�"�I��
����i��	h R�&��Iֈk�~aw����4�}����f�}�Z6���0��e���*#����Ce}y%��T(��4�P�o������YB�S�ѻu2�z2u����b�}-�g~�H(���y�R�]>K� Ƴm�L|��
�������6�xel1
�xG����7��a���c�
+߹�T�g��p�!�XP��LAG��ɡ{g��U�3��ᓪWsEl�6���7�&��>�ǹ�v�;w�nS�#;U$���7]������n��$D��aQ���s5����	*�Uxn���j���6ey�����Vz�P��c6��t$��+�D�F����*��:l���:���ʭ��Ka�-�Thm��K<���,H4���F�z�`�$�?e�	;��*7E�4;1ʇ�_��k:W�ob�9�B˔b'�|)�m�Wj�'�*;�q�}wE���V~\�ԗ	-��ۼ����!~oP�J��F�}��A5 ��h$;�����2����[>��؇zȵ�2���Z�Kz���:���/y*x�K>C��2�zJ�]���q��&-�W�2�UO�덦S�8���r�pe��S����0�*JU�6��P�v. �Bt�jު#�)�<��;��&�S0��C�G�����!�4_u�����������N�����g�A�0 *��ٕ��h�Aa�`D=��W��n�wi����IR\t@�I7�Yހ6#�@�C��Uy&��Ks_0�\)�h*	X1Odt���F۪}Q�%JG
Ȋ����L!�7k^�v�mŁO�l�S�Mn=鯼��y�C����̠44�q`�������3�8����Ug��ie�h�/Iz����h�V�4����A��,kRa�?՝�k�1GB�M
�@�9�����0���Qh���{~�@g���褨ngp6.��q��*~�?�oB�:�x�g�G��1B ��E�<=�|�4�\��ޭ�?n��N�O�
\	V���l�-�/2+`�{�+·��D4Ar��埫���9�u�w Zp3���K�{���c-��h�=�I�� _�H��ΐ�="�Y�7QE���S��7�\j�i�I1�[���GP��-�����P8�@�a�Ο�J�������uK�S�N��U��[oF�=e(,�Y�j�*�`I�k�lrk�<ê��f8�Dy�T��6�U<G�K�,�P!���e�5wJ]�����KK��WHz��A���u��l��*�vy"1#QvVm�bq���:��]��TC	�2�!�jn��W0��?��y^����	�O�m��9H#_�!o)��(��ۻ��#��F� }�ʤ��oZ�=�0v2�,�U$��=Q����[�I����ޤ �l�(ȃb4��^�%��ωK�h����~e��t�D�}F���(��3�:�s��tx����9�řߢm<���W�N�f��~ 
P�U7�#P}����z�����b%��3|�����ڥ��v����-�����>}�0�(+�%}q�:()�����ny1f�؍#k.��	?��^x�$
@�ܖt`�:��A��x0\�8֢\<���܉��}� ��?�CUU�A����'�1�J�E?BQ�S)�,�Ʈ���1ឰ��P��p��j��W�-����Л>
�B�|�"����G��󍂸�(��$�'����.�;��jF�m���S����cKH�c�|+~L�~���X���y+7��0k��&=���eJ~lI<����Xp焛-�o��8�G@l�{v��D��Ÿ#��ҫ;��?mr��ą�h1׎'P�b�#Ȱ�$ Y_��h�C�oQ�[� 
��}�ǉITK�R�ػkӺ��P�:ܚ����Y�����ĺ�e��[����t��#��E�!5
Ђ�q��^��q�{	�
Q��/�ci�9�?��:��z�_���}{�NNe�o�
 ]6��n�ېR#=���Rk�����J!G:-�]Z_D�r�T�X��ZS��t�������_��8���[p��ͽ�Ԅ��ԳZ�ة��ӣt�۫k�}��['Ji���6�R�л��#8$��c����h��1�t<�,)��9W�q� ����o~�Џ��z�^�[���:s����E�]��J�R\|��+Դ~���t.brCxb�b�v���"�+YQ��)�t�#(PY���
�6����i~7�/ {")wڎDG[�7Y����>k�f��>h�ԏ�[<<��:wO�g(�$a����3�%�5 ���Oz�q������A��쫪�
�9���L��4����^�{��j�xG�	m,�XF��M%��d,O����ا,թ�kJWE��mW���+P�ɶ�1�e1Xɨ5@	�Ly�C�]�~ֲ��\�_��o*Z�@�L��_Q̔XQ�t��J fV�3����@�/�{��K�?]6�?�]��a%���V��M\(	O��� O��Gx�1��E2`b2�{���H�R;Zqʤ�X�7��`0���u̇L�PUG2�0�I����x�EM",�G���MK�����8�osG����";��
!Z3~��eh��c������vf>V?�-c��R��z�� �2�W&�����f�Z�ӂ��1��L��u�32������Hjj�|c%0�kE�iqw+�UtT�u��|�����%��`.P�?�.�J�FT)�_�j ���!��N@��
��\p�,7��Za2�� �\EM�N��w���m/\��8��=��N_l��a���^4��U=�w�_.'P#xTm�^�pY�'n��6�{,َ��p�_˖ABnx�}�XEΏ�Y �@�T���̪$�-�*�ex�N��6S��'ɒg��`�&�Ƞ~+.���B�S�m�ˮ�]�m����h~�Ye|$��Y�~sK-��;���a��3NZ܁�UM�(o3O�3)R3tҌ�Uw�{� (�	2 �͓2wێaaqpR�d6��	�T�@5�CC\����?~���g���2��m�Bw�G,ҭ���h&ŰH����j��J��{O6$s�|�.����r\�Q�w�#�3���5�U�KH�����o��Ud}�U��n��N�4��%��L�l�Ŕ�6ۦ�?��P<��ycdYdt�U<
�۷�áު�3Wd	��bk�t���UT:@4%f�(�W%�A���)[�i�	J�C�k��qcj�!�E��I�aѶ,��#�h�Me�H#�
�8��9"�4xg�<���;v��M�v�GlL3d^shh��s��vjzb��/���y?�A�}'�����N%��?+wj�IdsV8��TH�1�פ:<I�]�������>k|D����m��e<Z�/�[��9��҄˶�ٱ�w�*rTIi��y�����q�0�)�e��k�����w�T��������3��u@m\o[����A�y�����N�;B=��vP?������o�F��\�Ro��ⴚB�a���P�j�������v�g�i�-�.ʚQ�\k1���������̇&�8y���ZS�t�3�7��V@8���Ez��L�y��e�~L՞�њ�lح���z|.Dˬ/���x�e����8jY4�Me�����a��O���L>E�`?�°K=���8�A�B~�l�n?b��yd'�Bw�*�u�w{�9YB����Nʴ`�N��P�����s��z�#��B��E�pϲ�\���n<�CyR�*7X+� F�8gL"V����^_�i��CZ�*��O��8�.��F�B���xձ���+O��4G5��І�dlޡ�W�3\[+��v��z%�� ���'��\G)�m�9��y(|�M�S3���8%�� ;��x��}5"Omd�b)�P0���T�GR�a���H�F3��Q*]�]'G���|�Q��%<L���%I�y�D��%�0��v���=%[��?�c�%�}D["\���@uB��1PL*���]�	��=n��nyf���$,� ��� ����@d+�2�U�q�.����\C?)��j��V�"]xi�x�biL�*O�E�s��u
;�X 	՚�.�����A��K��!egNZ(�Hv̓[Seh����?#�M�Ƹ��D��$��Զ�xm#HFƞ�XgV�6�=�DA���G?a]*�T�s�[_|��:�R�~?�q�M�#��N��ە��Lq���ja��h�Odd��WNaYfo�L�XwT����1✰XΞB@�ȭ�ρ�6�&Q��G�i=�dk[X�,��껈F�7�ŀ�i�p,rR�5��G���te�seP,r�ƍ�����Q�7޾^�0����-c��*z�O�������q/"4�0|���h:��eW�,߂OZ.h�B�rg�z�n�z<;:������Q�Z;��<ݰ�,�)ؓmL�a��a6��s�3�P��ɢ``r�zQ#D/��Z_��t�m�c*�-J�>�õ�=�vu�>j������Ó03�}!��4p�"�6�'9X�Ĵ�]��Ȩ�aj��E�uK�H��sG{�D
!C�vw�aW���@K����{�y �]E��l�A�w����%*�n�T�{��@������2[V)o�|�?���]=6�Hn���<��Rr��M��t1��pe{��?�e�D�\ݧ�;=1r�쑥�5[p{��~�k�|�w+I�4r��M�!�	�.C�n�ł*���M��W��s`�
-����s�6���A��S�=5�ON�1X<,�`
]��C���̽���(I�'I��Mx�]��ٛ1F2���gh�_}��q,�+J��R��:�+���U����Yy	K���F
�'�Ɋ�aђ�Z�c�F�N�e+'�8S�r	��^��I�A_��c�E�A��������)�PKŖP6���}�ӽ��a�zO^d���A��SȀ��F���o����lV�!�I�ƭb��߰w��g� $�`�h��d'�s xϕ��Ɋ�H�$��ӄ����mk�Ń�Yg_��+�ڮ����ͳ��G;*$���l�����;����gy`�:�N����И�!�$��YQ���JW��$`��EeW'�0qj��i��\$;j"jl�����NI��C��.P�x��:X��g-��h�I��P"2cF�Kg~&��à�u�N��K\��7Ǚ
�{"\���e�E�!�U��]�:�L��M��u�@B��π��VS zՕ�'��96^3�".;�ICvF;Z��q�g2'Dc���φ�+h�B�����#3rno{
K2|�p ��#t�+��u���1#�S�H2�ye�f��t��ɕs[p�A4A���Wp=C�cWyP0��v�\&�Νfu��g��Φ�Q#{h(`5ImmA����X��F?�J�2�_��"&��ᷚx�b������`ft�o��[JQ��[!�3�)x��B5���ć�$�y)��n���y��D���u�0�>��@�������^f�dvٴ�x[���ّ�h���*0𖈼`�
T�;NДpqmH>̫�>�v�5�cݷN��V6:&ly��tV�~~���AK	�\��%Q��g!�E����K8Eksp*�Է�Qcx�ikE�ݤ	��2��'M�l�H���\YI�����-��kG!����)���!�C���FW�o��֖5=��bk^6���g�P��}����ϲ��|�o�:�-���#`�S���(� ǲ�ء�z�>�Q�-���+�3`e�^^�*�-w����v�U���s���BH�A�⤊�c��+!�[(I2s���I�<����q[�k�Kg�YR˙���GM���#� �c�k�R0�1}w���A�K�!3��ޚ��xop��(Im]T��Oh|��#D{Z�c��u>���T��u瀛��j�!a���)��R���sZj� $T���31��X
����|o�PO2l�P9�Ĉ$vb���F̈́�?�4�2`����i��;�b2����-�ec�bI��?����p8�V��Ta�C��ⴸ����~?��b��h�� �����jT!m@YS-�Z)?���h�tV	��J���P&��=y�v�?�:�'��2���
u�?<�vKOШ��dd��|7�9��,�SŎ��ع�1ɗ`�>���h���m|�����y+�Y:�0��q�9��`�jm�4O�8<:J'�����+�dqEBh-���ۇ{G�jO�&���l�d.0�!
-�=s?�47�x p�y��B���X����ˬD]��sAL�~�A�Ǎ�X��?3Ȏ����3APG$Z =�TJp�l&�a���&G[�yJl����$q�ᶳz�3���[Et[���m�t��Z�Oq�t����O��ӬJG������� �oƄݔWk��0�������dr*�J�=��;�dxs'=z�O��oddi�'�k$�GJĈ����/��;�7	�\�]0�ꑿ0r��z�SmR����b�@>�����"K��DXQ��gE]�����I ��.���W�<2.�wV �B�&�F���ss���������u�#6�Erf��)CK�4������h{6�
i%VOz��D	�Y��x��X돂B��U���5�����¯�PJ��(iz5_� ��cך'���ޱ�� �����#=V��
�l�³ ����?P�~|}�S�p��vk��t���\�- 2BI:��m���!`~�2B�8X��xC�|�G���O&�i��u�[5�Y�0�H�3�y�bv�����(Xff�*����}��r��iQ41�BhR�B5�rm%���g������q�U���X�D��07�>�IW�ΓC8иl_��~�̊�caZL���\M�c�I���U�́44�So!�]c_n�+�������� 檂':Hpu�C�(�U��ۅ�-�{!CƟ������`���w����;�oe�:o-�E�3�y3uF�E�s��એ"�Ű�n7�dߒgD�*������f��}ǆĩ�$�|�r��t#�H�� �1Κ3�ԯ����	l"9(�׀�q !��+7$9�W�rK�K�ok}f�ND�R;�Wd��#��L�G$�%o}�b�SOۤ^�-q�53	6|�T[����@^�n��o�Q�����:�%O�C�9$v���7��C
��h�3/������wŢ�Z�x��W0R> �bL��gt�����vp+�+�*Q�_6�2w��8;�� 7�i����:���GqyR�U"�h Hss'�$	_���6s���e5�i4q��B�Ď%ĳ��8�/n�܄ǧct��0,Sm5p��A���s����� ���w��=E�S��K�Q@�����Y����k���~>��&NF�8��#~�Q�������5rF�2!��^)�����/��Жz�%����^��DF��}s=��G`��������R�G�h6���(��u������p�hq/g��P����&�v.�������S{�s�Ab��o?��-�R^�Y�8e���%*�f(���;8����Yڼ?g�:��i�ℳ�M�-�P���� ͍��6짿;���l�Ubf��J�º�0U׼9�(jAWu��������e�ь&�W�l1Ͱw~�r\�-XX�c���GTle�mF<f��-�	 �:�/�q�}㤽�{�tr�B���o��~�r�!룻|�7��s�XW��%@=y����o2f�hhE7�P۔R��m�q%�{� �v��z`��(�u�. ���{�V:� ǇA��׎L�߶���Gg�;	8������g�W#{���e����U�̤ZN��L4�����i�NՂ:h�^f�ΨF�wS3�FM��S�q��� �y�P�J��������O-h��^�]h��^l�P8 Ta�������f�Kj	D��J`�pJk�8ǃ;}4�k��+ߓ�i�
w�;���HZN�r�����x.%�ɗ}�&���J�/�Wk�I���~<DK�dcQ��~�3=��A!�p��9;h�7��;q��?��/Zѹ2;�m0cB�s��u�՛`ݱf1-� x���G���L���t�<����\����ay�V]�E˰{�d��)k��
�c`�PJ�o+���Ms�G�� U���N�]+G�Y��А�T/���M�:;�7O�{�GB.&�D�\��d��C��3�c��qꓗl<������X� o��p����#��d�YV�UZzi.P����T���S�ݨL�Ql"�y>�|��`��K��@6@��q9V[�A�e}?g�#��~���0Xt�<ϯ����7�B]Bݸ2����a�%�PD�'�W��<X?J�/�yG��~������.[�O�}&�M�vj�/{$�o�@l[�$y���f�nm��\����p�BXzy^�����������)�A���	��$�=���n`m�=��w���&��홲Q�璓�m9�f.pt?x��	T����*,�!L�u���f�y�eƭڜ������=�5����NC�� ^�%
-σD�\k�y�Dr�Q�+�H�� �
`0@1�e'M�6$����ѷ�	��P�I"��yȨ�p׉ω��F-{1���,܊ј���z�?��#h��o�0 9���m���~�q�ջWc��F���	)W5#�6/�Mu�}�0�H� ;S]��c'�\�!dt,}�qv���txTڣzCk����ˈs�BF�'"�S&��%"Ė�R�ئ3sw��k�A�P��k2e��?po�ټ<�KiB����Ҹy�@D��j�7�T�WP�d>SCz�o��W��z�;��'Է���iyk��*:�)����}�=�� ��y�M����%�ѐ��担R�,��Y䝋D���)��:/�s��*6���)8�Cꁬط�EZu��Q ��2��_U@2�|��f�ё�,H��n��%%��#F�ov���6��w*ץ9����%f0vY!	�ij�$���w�	�6ʮ��_G�wΙ�=�¬,ѧ�\�!vԪ��_����.��)�/z�d��!��B��o��ٛ��%�r�J�/���/g�KEˬucb3¢Jy�=
��U�0�V�YB��v$�n:CAf�������m�o"%�C� �7��W��mt��������wFHa�h.5X(����D�j%L�5�h�jh����G�F�4������}�4���.���xWe�b�]�v�����o����j6����R{�'O����,�L��§�b�$+��_'�Z�H�OMJ� c*���Cd��@x�	G�F���� ���S���&�0o�R�pjXioż�x��V�UqngHJ�*H�Zh���"�*���~��u���v-���f����V���N���|Q�e�ۥ�L7���.Z]�Zt���a%	Y�RE�K������̮㥭���a��|�,w��O��k�2>��a8zH�/�>܊�q{^D�S'�-<��z���O����������k|��So����|�WrA=�*
P^���&�I J��\�m�zO�4��7H�N��"�����.(6����v+�����kn��+�e����)��8�J������{�2%e�¼ݑ�h��j~�؅��0tgbۘ-��0H��oZ%�d���*��$k#��ښ�G5��!2������?´�me�Z̚(
	��I�t��m��cY�F�c��à��@ܢ�#uډ��׎X�^�Tb 0�l���{k��as��{�5�yD �i+��5�E�cŔ�� ��[ob���������	�s���b���Ur�T����F��S=$.h�9������Y
@BBǆ�{�����e�:ɬ��'�l�z|��ꠛn&���R�hb�)X7-9m�7j��%(H
�'�9���p� �"�}p�s�L �eek%{,4+b9�Q ڬ�~r���#4Uo1��B�:\w�G�"%�cj��R���'�r���D]���"_���P��WD��L���N�ݦ�3Y����}9o�x@wJ�ʭ���<d�z �����_�McۉS���E3D}��n�X�����R�ӊpJ�
D�8� f`��J;쫈�Le�}Q_A�(j0,=N���-jcL΍O����}�ݤ����󾜛��K����=����̜��CW���3rJ����[�����*�RA>w��b�����^3݉�=��}��ZEUb(�a��.����-
�7�����4۞�b~̫�&o;�X|f��������@iΉ(ݻ-~���6�l���P�s�7��Ed�z�M�o~?��r�����a�F45��D�)x��דXq$4&h��{e��at3�k�; ���g	P�s{�6�Q G�0
~���l6P��կ����t�/�����5O�6��m�Q��@)K��.�F��r�o�'��C �1��N]*/���c-���BI� �_�x�V�=��,֓��������kE��I{�WoDc��(-4L�?:��`�����:�Tc1.�Y
����û�A��tw�x�0�}��q�b:h3%��_����3��z�+����C��"[R�)��k�B� UZL��>�"l9�,Q�c�k�/巙Pq���h�q��w�g3H��o���E˩'�$�EF"�)*�&k9k�[�k��zo��'�s�Uc�R*y���v�$�ۉ�fZ�ݎ��!����+Vt����3hcKV��O���	/첮qE�U�
�JQ��*�E�Op`Z����>���eW�k�0��a�T�<�W�m܈\K����{�� >����a$�	����MqJĹ�
�r��n��,���B�r���#Ȁ���>M/׼��r*��/Z{�V�I����N��0����z�u��\����J��<t2О�`�ǀ�W�0����2�O�ܓ��A�g}� N+*�]\f<&9�%�4�l�����dG?s�{$3ނ�}]�JW�Y �~��^l��_UJ)�_cz3b#Rtc�l�P��|4$���8��#���IU��N,fP5�mc�ǧ]��c?[��0
�(W�(�D�֠&l����0^�HW��i,�R��!H�\p+��r�)~�H� �D}���۸���-3i4�#�[�\�3t��'��&VJ�*f�_�^�y�e�۵R�lZ���f�r ���{�J��C6_���zj%�G]LS[a�L�>U�"�L�c�d�_�Gʎ����#*�7RA�zQea��֣� �H��*l�;�t?ֹ��ڮf��0'�+A�&�/L�p�9�Rc�i���*A�-z_�i
�샛�Y�>u�]��F>��)�O~H�~i,���L�h/dC��n��@ 1�&ȗ�/5�|(�� ?@�%�S��D+h�x���ɝ�]�߄�3+lK�oT����Й�����ވ*��SO�=3�nSe�S��N�����&] �\/ch�,t�z��!5�I˞/�B���S]�wO9X�}AJӜJ���Xw��JhY�M���)���(����43���	z���_��2�l8;���F�7�o�X�W�K<9��!��)fa��������!��cK���d�t������G�@qx3D4�y�F�E���¤���K�HA������0���ӎb��?�#K�=c&	@�s`-}��CFgY=���\�ϰ�Y�kUFL�;A�%��"3+�p�wH��\Vmf��e�bSL����!�<=3I�.�7l�Z��\�����)�>Wo���$푷ЬY	���M�^��	�SN�n ���f�3���O�J�w��+�?_PTl�?��NǠ�������M��Z^\�#J呋�km�<$>�`���W�=���}B�ik`���ݗ�f��U�o����!M��XA<�@1M�
�{�ؗ4�H&~LzC[�
�e�22O	t�>`���ѣhf!p�>�"R��� ��aЉqk��ꀇ� F͆�MƉ��� X;���9�TU(��h�p�M���?���S�D�rQi���b!Kń��^�^��t�HLĀ��N���	�Zi��aK�.��G����Zw��`7ŗd�m˨G<�m9�}�[���'n�A+��VYa�+f�-焽�k<C_����,��$_����[f����Yމ�[$O+�Ĵv����d*�l��-�pgb"Ԁ��v�3��v�֛�P!}�X��,~������3bǐWja��t|c)F���a6�������'3�duU�f���|�E~�FV��)�{7?m��)y�O�<�๬�Veѓ�.Mb����"P�:��Б�&4v�H������n;�mҚU#���r�Ց\a�J!Ri�R˖��A�����B��/<�%�I2�eSn8����C����_7��HB�7�?�j!���3�E ����t���C����4�ՁR��gIJ�׿ ����FhXv��t�3�ѯecEFl[�q��V�<�d94���|��D�4p��Ѡ��s���tĞ3��Y���/w����W�d���U��'H��6�%�?��/��J<2�}p�3|��%.7�\�XZ�2�O�1��/'7�NmȒכ��v���%���(��N�"�Kj�-ZN�y���H�������u�T�ӂ���V�H~�H���EG����fv�!���g���P�C�1{gw���os�Tw�J��_�O����'>/@(�i9qf׎��PA��8Ng����`��A7?0n����'ߟ�S�M2���^��FcQ2�eeT�p��W2�F1�f>3���$Ņ�l}�{^ zm�T��v���۫!=�\�����F���ǔ��$-���s3�|F�+<�
ՠ�8s�q�1Y	6� �&T��5��*3_x]�@� ꒪��d�7:�U\����D�\���>t+�н�B.nw��:��׾?5}�^]�KE�FdP�jWK��z)W�5�!���V���|�KRN����������z)j�.,@�.�*�23F�/�r⁰I󼈷���@�TR�@L�hM����!VP���a`@�s�FB�Iw	a֣͢g𳥟����ɺ5|>�4q��/)4q��Tsl�b�ˆ�U�U,�ڴ��.F���Rt���?�7�2q��L���r��7�\L7�DG��#���xj>�E����ͭ�hP���k�0ʹ=6ߢ�_���i�}m�.?x�󧩥��KC��Ip78�K�~�S)`�(K`������yW^�3R<v��gr���,��@g�@<]�Z>�(���'�gBl]����m��ݥD��ʋ��E6N��?���Rw���5y5ֈ�8O��(�Xܡ��"��Fh�C��-�u�X���W���[�q߻��+�K���������lg�$�gl��4L5�f!~�k���}���e�.t�K9Δïa��'�&��p�w���N�΋U���hv[{��k�j	�Vn�9�G��EᏫ�u;vv���i
tr\,��G�L�t(y�Fr�(����t�[0�!x�V�RC�d�w��6��(�G��\�����gAh�4X�/b�g
��[�[@�n����`cf��d�͢�O����;��.*��}����f�l�K�fA@���w?x"k.A1-vz�s��*%���S��͟?��IJJ����z��[�2۴pW&�G[gS1�M�:!E������������6�
�R����@E�dAOt�C}0��:*5�Y����Z	h�(��W�yg*�m�w�k�$������!�oy�i�!qC6/�6*Aꡣ��A��A{ۤp��g�䨟�~����"�Z>a�LR�y �Нş2�-x�qt���߬�-���u(�z�j��G!~sx{��_^���[)+�㧥���,"�er��C�gV>�'�ه�ţsa�^=�~�c���`�x�>�dX~媤V��ѠM>!&k�wH;��P�f+ ��g+
���;�U�j+KʂS�'[׈*آ[ϰ�k�q��F���Í6/+�\� 2�ɻ�5 R�d	�~��V�}9:�at�<��C<1�v=D�
Oٛ?P��V%xG��$a�� U!��I��/�6Ũ�u:����%�ʝn���'N��a%�D�pݩ>���)*~�@�}d�8��.���W�8vЅ�h�����Ŝ�6��7��d�̠kA+sC���l"���<��1V���%��(�FD�,C�F�#������,~ۥ��^>���-rv�K����R%ϙg{���s�$�l{���ȥ���<n�gP�Ru�����4�Nɢ,yMa{����n�H�˗��p��k���:л�oj(�D9�?mQ�ْ�%7~ՋMjK4]?�v�4���'����ؾSo�Z��_�ch�*����y��RJ�d_?�|Rgj��꤁�3Xp�s O\�{A���!}-al7���1�=m���]�F:S���������I�PN�Ý����N�'�^(�KLC�#�2s(���6�9����:d�O⇞b��No�m��|�*ô��-��H9���N�9Z]��lS;Lb�I�zJ�5ח�}�Q��d�ЅK;�~�X.�O�NuH��2��R �ۿ��1��1�IHׅ�����X��c)
p����g�)����L��(�4�$�j�IvBړBfӶ��D�:��G���3G?b%Z<�]��2=��@,&a�Y �B��[S���`,�H�'��"���-�7R@	+t[�r7�`�[��Mb�ˎh��*��cT�2�?�1�mݖB�jQ� >�䫇M}�����]�QD�l�vQ�ѩy�zT����~�D�p8�AK��C�1:!��g�����W�{��;)���&��tO��-���hd[F5�7�<E�~`��{���o�z	�CC���-q�+t��'�Jg%�׏�rk�_;��������GG�W��Çq���۹4�<GFn�]�)��q�lp�����6o-٤�"����->ЪK���K�Ԫl��Fa�z�)��%(%��+L��Εܱ��h���I���S'��HT+� �ɖ���{���X�"^4���axLB�#�f�98)x�q�"��������J!������t鄿b/3�?q�m!t-4[���;a�v����]i˼�7��݆�轋45�F}(�`1��Ĺ&Q(I
"��ە[�!�$�\�I$z��.�
�2;W��� ��L)��7s������=��� ��?REx�@�����7C�<�PD8*���ѝ�]�; ����A��Aw��#�aBvg��{S�{���ڬ�v��80x���;,��GQ:TPe�yN����$�_�� �C>5i��4~p*��-�^r�|.��R��'3<~0t����̺��7"�ʄB� ��ߔ�`�����ڂ�">>;f�2oH�I;���d�o�E��TT�&O�4c� ��o�������]	��2��@�˲�m��`���ZM�����a�Ʊ�J�t 1���r�$@p��������/T�^�)�=2���(7Q��M�^͉#�#t�J� {�|�auWv�^�G�g�B�èǁ�n(l^I;AS)"T�bl2겡�[�O�
���=A���fo���T�7 �)�z��`���3۹��Y�2s��Ta�b��#;���mO4\B�6���4Ń�[�l�-�[�zM��ꤏ�9��)�r1�v���c��V5ٚ��&P��T��Vw�ŝ�O��D>v1ډ�4��R\�~ ��h�Ҡ�/Ǟ�,���Q(d����Dd#UR�T����M��̻��#<�N9�Z �~н\����_z!�o�@�/�4!�Z����k�����(�T���'�B��tͲ��=/�oX�8lv��ْ����S8���6ӣ�_l��j��24��>3�@~�L�	�$f?h�.4���+$�9��W�	le⿴��=[ƌ����>a�W,��v&��
5�{�v������ϻ��;5�$ܐ��6	�Dv�ېŬ���0~%ֿ7��Bp�����DW6?���\���>��B�M��7���SJ$k:Vr<��M�v�8o�2��U@�����!�١:��
p͔:iQj�L���-��o���؇���pr�>7�����	�� @K���xG;���֚�G�<�\��U:?2$<��oI&���p�{1$BA��������4����^�,v��Z|�bf���3�!"���cQU]7���2�5�dW7�&��GE���g�QƧ�1������<�A?x���[T9�|��7*ɑ�p�J�=7�  �\���oFh' �#__��䧨mT��K�Ξ`Y�Գ!`�6�y�4����y���糍і�0H%l(�T�����Ɨ^� �l��%�`Ý}'#\"�W6Z6�9�}�C�x��eq�K�����n��]-)C��Z����)���_�zO��^i�U"���4���2�G�l��=.��ڻY��P{��e]]7�@�����C��Tq[Y��vԶ墤ʮ���F,b�������/��i0���OUM>����[������WN��{Am��C���G@*'��G�;�g���{�N��~"�v����<�eK�{_@�<�R��\�=5��\�g�t�Y
�>J3��)e�"?�:��  RF���]��k�����?���滋�i����x�pB���߳~Vo���o�GT��ڤ�:���T$P3�����Q�k��CȢ3ढ�JX!|�"�G�i8��XI�:�'��.�u�4	ɡ�9���qe9
��a��u��P�Y��YT�EQ�,|���?E��f=O�~�Hw�'
%C�Enku9�#]�$,Ehs�����~0=��Mˈ0�Y�Y�]�s*�6��x�g�[;�OY�������E#B*��a M�F5�ԋ��M3l���p%�ķo��Pd��z�ZAKX�B�@�%%��A�*���b!l��{0%�?���d\j�z��u�/E�9x��N��	(�kb{6����h�U�e5K}T���.�ј���1��� �M��u�W�Q�M	&��殂�Ю��@4�Oa�=`�d8������g&d��$��Y�C�!�!W�� ��*��r05!���V�!��N0��X�)�m�|1��4��ݲ�S����B0@��/5�L{ƈ|v�� �С^����}��2��^Re�q�Z�Ѕ#���_���X���(��:����<\��������{!���m�S\�U��2Gd�_�
��B�՛��Ā30[5Hki�i6���n�
=j�){�V{p�.����#<�V؜�#��Ra 3X:�6���fhdyr�Sy�%���xO?��ޥ�渚�5�e�J��׳!��s�(�pz��.[g�O�����G�X&���1u�����yـzIY���lP����$�:<��j���TK::Oq%������[zW2��(�dE7��a�#�+#�S.5}�3D���瓧zu�J>l����ij��;��� kѰIX�θ��N���8���r ��%!���zepB~��;Hؼ|�^
��0=o1��\�E�¡�{F/$h����!��?*�JY��B��PM�%��;S��ǲ���W�V!�>OS5�����\�_�7D�K���{�c���Ġ9�*]ԏ^��8�W�X\��>`I�]ܕ��>z���7��D?4㐋E�o!�K���Y���C�P�NwzQ��o�F�m�YI�!4� 06�KJ-�@�c��>Dvj�~6�H�V*b��7�ˌE#�D�~�����]d'�G0�Í/�0�e^��S6.��:�T���O�ZFP�h�C�g�Q�G��0X�>g(S���a�l��C� ��D)�(&B����0�d%�.�;*v�ϣ��$~�l��41�� Y�?�A�h��<A�;1�Z�M+.��n�̕��*zYb�g�zs~�@�p��N�u��:�{�@�-;�´P����n�{luˁ����e�1C	!Z�ug����M�\�<̋�Rh`�hAV(�#e·�D�_�1�ً�r:�J�l���Fr�����qR�p@��y�i0�-�к �����,=v�!��4�W�pYL�$�	M-����r�Wӳ+*��NW���u#�p�4�]���?V��(���&�z��a�4�mpZ�^��@d���Z���N֩E+7��6��#hYU��Vaߐ��%V�ŝnU�c���+�;J�<��� D�܊54�>#mR���p���,1 �هJ[��8�a|i0M�{L��%O`�Ժ�k�<���&�i�;��v�ł�;$ACX�(�M�w��#J�����jDk��׀$=�y�>z7-gs�1tq?w��R9�̹s�}cwB��:���F���)3?\G�v@ڛ�����^I�Chʠ���G6��S���7"�*_�1ZK� bö��oX�ix���77��;d��M�1��"�|ޫ�	�Q��L��A��]�p��U���'y�;K��H���`��+q����*2@�Du��j��{��\�"��� �jSD��>�Xny��*$w8��F�jv'ë*H�L�L*'��񅎨@`��k�:�Q�5��Q�p�{��[*����n���[~�.�p ��O�)6t���i���F�g|�r�X�0F�[�g)�4�N[a���ҝ*��#Y�$'��W�H�k�C��/�����}�j�lی����@���l��cTA]l�HYr!��Bo~������GdS ���+0��F�:D�bX�9� �����y��3t��:��(�;�g��7u'���탙�>��5�7w�|8�(��3j7y��s�Ruo۾YFpc#�3�=���L�;���jWK��
�%�>IެM��i{�f���\�b>�;"��ٲ�gS�!%<��)_�Z�*�R}���N'MH�Cx��*4B
&8��7�O�3$K�6�_���?_J`2q,�\p�����==�\iT�<-��L�pK8���X������_�G�Ex)?O��o.4kt���k\��O����,r��㯪��t��J�QE�@�3�:)j
'�Ͷj{vV� U}���^I�bV�)^~��ph��f��M,�>�S��t@��ֆޭ�8�|;p�,e���p�S�A�%���R���"d�=��N5��R;q*�`�n��U��ڍ@�(\;q��ѐ���`^�Ќ�XVf�UEG/�Q��7�u���������p����x�+4��s=Bhr�z��f�wk��+���i���H��h%���R��Et��2�7��t��-;"h���>m#-ڂ�jY��0�W�<�w�"y.��5w�"���;�Vߙp�8���W"�_��O���tA�@.���Y� Ve����X$��fuq��4r����k�đ��{+a�DH�_^`;�@GzwZ�)����iaͰ%��c<(��Z��Nqq����G�A�'W�li�ҟ�h�gc�`J�Z���S�tְt�x��J�u`gd������~=��:N�vY�}�Œ1�.�.]�2���a|�XI��{@�c�:U�U�'N�i0S�amT��橍Q��|0�g��y�K��aQ%���v�P����~{౔UKE���X����,DDT��< h��hFFP�<�	�f�vɤ1��T�0��|����h�3����x��:Q�,�1��^*���uKH���=Y/������ g�0�>OE��H6�� ��B�kz�Pl#:o,/p$X�|�����)�9s��������Ï� 'n�~&$�{�֐��39�E3bO���XĤ#��2{6+�PSBv�?�)@�\��Q���ݿ�����m�jUG8Q��t�r�C���k�ʉ�@{�\�֭G�S���~����m:��,R� �܅��ˁ���h�C�J��BT�obb��x��;%S�(�Ac↝O6"nfBD��5�|�LF)g�0Ty��`�JnV �H) ����@f�ſ�[�N
915 l�gJL�gQJ����y���A�`�8��D��N4�^빕Q�/�b�oOBJ�?	T�(/��HD ��z��W���]~��3��y�7�l��D��'4���������c1ŌPUy��uqz/V�J�Ϥ�]u�W*��!{����H"6n�fpwy8bF�2�fMF4O�bP�V�~�EP���|�{p�������/)�u:���xt@8�ͧ�<):ן����!�S�dzi�)���"� ,�h��[K��|�4q���6�88�|g^�[�tqj�����^���J��C�,)��c9^r/+0�K�K�]&)W��;��oCn� Ic�Җ��կ�f*�5ט*I(b�/�yi@i���������*��~��Iҧa��!E�}��:��R�S �&3��sK��	0�,��5�\[����H�^ԟ�{:F�����k����of���y����"��p����=1�1=碴���gV�/�4� ��m��۳�~���|�:N�"0�T���������̋%s
]ސk��1�7��!�O����x��9��7c6�����n@�u�;��	�)g�*�v_�u�i�z�P&ڐ��0� �r�h����:߾��Q�y47��� f��蘸�R���Ƌ	G��~ƈ�ᱰ
ctUo��(y� w����Zɢ&�VJ�=�^����=҈Ѣ�I#�c▅Đ��吙�?v+E�+�)U��-�:�n;���>�㍉�ΉJv�]
1/�SKeإl��皁���F:��m�X�7���7!�nu��������p��C�� ?�j�$N� hJd���Nv�?D���p{?�'\��2w>�'&�8į��ս5��u7m���3��hX���X2�_�H�5�u�)�$��P�?u���L�L��:|�x�����Jg�E8�e�I�<vm 旋Gp�K���!�IhM[ہ�ٴV8�]��?� �+hՠE�i��k�������_\��
[{U���$����~�7q*\��V&��/�-a�;��Aޭ´���J�1A���,��աaT�y�)z�9wݘ���-#YM��: +k ��л�Z�|�7��Iyc�v�L=D��ݩS%U���tٿS��\��Ɛ��4KD�WX�S6�J2��fPb9��>�m�4>O03����b�M5�T�Q�Lr����L�Mʼו|�f6���g�+����\���^�w"�]�G�?8e{T�Zd�T}�	�
#�mrhU���&��A����ؼ�6�nF^\L����&�Z^dA��|�~פt�#�d�i��������"��Uж��5��>w�q�,+�����ܥ���z�oԤ�u��
�=j<�BZ�BU0�y'9��nb�{~L�9��<l�[#M,tk<�����꜑U����t#_{���
�w�j���b��$�:+O�a����C1R9A�ĕ�LK�YKn�-N���V�����DI�t��c �U"�_Z6�)Q6��-ɞ��B�,L�[�2"4�5.�6'W��`������}�,K�ͬ�����G�7|K�1v�1R�$�fVB����k�4�5�/(��c=�42E͇���ʎV_���
µ�ĩ}" p�B)К)�l���X�7������"��u��-QڼQ܏U�	�u�u:�V%[*_�C̈́F��\���^E��/���;�[�>��)���'�hT������X�{Ѽ-����yt�a��1��"���Еiy��D��A��h�0��2�t�$��S[ǒ{W�ޡ\���c�j�8j�,`iMY�)w�����]����fq�ݷ��:�ܩȪ%4ɒ��ꨯ��j[<N�,�k��%��VIU��>�������1$���= I]ny`����yW�	�F�#q@��bո��Jo ��G(�+ΤK�o�ȿ�����iɇB�5G� ���ſ0�H��f��,SE�n;�Sg��qq��v�߯�����Ȏ�V�|?ޔ��{��04ߙ�e��������g�EV� V[m��^}KLED~�g1W���Zd�8B���5T�q���=A����ܯ��/��m���&���lY�E���	�5-�]'!�O$!w �P���h����B��m��V|e��<����{�H��W;g�B���lOz�x�_���k���3J4�.j\Z�{SљrW\ծ6E�w��9��xK�ܭP��-.Z-V������4�;�ܪ�݊���ԙ�I*N`z�)g���=������P�y��,�В���N�>-L]	�M�C/>�<d�RwpLc��E#�CC�
��GG��x*d���}K����<^<�
ү�S�?��R߂p��j�����_;���?Pf�5,ײ�Cޛf���2lAr�%�J�[��)lB僄��K��Ÿ�H�j^����|���tW�����HzU[[����b��t������j�v�Lcf�+�ys[vy=	 z��`c jK,w�����&�v��������.#��|�x-̎�<��Dl�ߵ�& ��wh�Z--��>~�y
 ,��Cz��Agv��R�@��R��m����oד�^|�Н�|��F�����{���<��A9�eeD��5�7�溢�tO���e��k}R"�6BT����
C�1��=�Ҧ0n��ɋ0{3Yc�cz���zG��5�A�2twHӑ�ڄ�0nX��;�=�v�������*�h�ؖ5�"#�މ�Ł
��`���
��m�t��C�k�*,���K��j7@{tq����Ά�t���ݾV-��9�vyzx��ƚ�q��6x����^f+��,�J��_M%ˊ� "�g�_�({����B�Ra3N`��P���!9�D��&K[:��Z�B��0�G�����3B���!'@	%@k�"\?�隲k�΅}:���lu���eg�T����9�a�7��q�ac����u�񢤄(���,�(���`kE�#�3�2$ݩ�W���4�-=B��	��l���+�h%=�R���T��Ԑ��|�LG�����?,�$:0a����Q�%�#�zϩ\iX�
��1�ߐB'<;#3O�wwt��t.�f�"����'�J�`Y�C�Kc�^��G�Jd����	dy�~N��������q�P>I�}�H�/�o?�U-׀�Q}<I������V@�����
q^e�oEBn�j��$���&�g�;;Mm��fe-i�[r��zSv)����x���fꪌ�����9��+�`�rr�{�WƊIؔ5�.9Ȟ9�����S(���Ԃw�^��� ���9��k��E�K�;�f\x��Їuģ��6 ��~I�*/4;��
����c)N,�d�:�?��9��}Lo����:K�'��s��x
� �o�4�Nއ�=m^��D5����� [�������I�IA�I��(-?�, �ɄO[��ZoW��"}�ʤ<j�\}>j'մ��������>��[�8���0.*����=��l%�N6��/����A]�0���D
�0�6�΁�Dwۢq�c-��d_���}i�1�����fG�QH~���f��+�@_�0�Ԩe���v��ԉ�i&1Ɉ�nѝtk��$h���R4��`Ɏ��l�wJ7]���!���ZU�@B\R�r����>�����<�난J��G#�f
�� pZ��w�����x񊒑�Yh�"_
y��Ί�k~;�A?���cO�j{wsS��3q:�[㌴M,9wvBjP�,��߳��9�Q2Z:�/�c�t���@�֬�G�$��I��+<r	2~2)�6N�;��7����S;I� �Nt�V�L݅	���'/��;�|-T
���з��W�*��_&�kW�F�,%�Z��WQ?� �ǀ
҇s����7�gg{}��Z3�o����Y��F�	{st��[�׷i�^�4k"EOڎ�����l<sͧ%�b�1սcS蹛������΅'�r� �32�q.�5.�7�)� �6±� \�ԞEA\�FhV��;"�ƫ� JI�GD����?����Q���IT���e���_�l���b��˱9j �(޼ګ�*U"��GL����Ic��M=ԌW��eWQ�IL�"aVe�P�ʋS�,�X�ca 7$��1Д:/������WY������� ��/3����!oor�)��s��jL4i���	���#uI���;i9����ʨ8e>|������Z8F
9����3��|�����ҟ�#����j�mk%�ᄉ����3�F�%e�20	�l�ݍ���ȧ�HH��t�QY(�T��4U�c@l�.�	#w1���@=�]+��B�k�6�!hOl�ߢ	x��͵��CB�f��g��=���)��#x�����$�/��4��%\_B�Ia�������v|�-X�c?�e���ZF����1J�O��W�7����!fI�'�m����EݖN��h���l�f�p�w��\mEZ� :�(�4D���x���*�ж�b\��E�����{���)��ZR��-�ޯM��;Y��PvN�k�lwp9��?P�	�ڋ�<	]�lާ��E5]04�Xa�JW7��P���C�H=��+����,Q�)-'r�*�����tr�)��J2P�ʥ\7�il������i�t�E �W��EG��y	�78iȆgp��MK�,��
�?_vgY�*@�L�[	���g�)7BЛ�� �>	���cB��:�v�U��j�P��<�L�)�e���<6��Tq}����{(|��MKc�
K�����=p��4~62)�3�@������ˁK�!��y�ZD�ԅ�6բ0Дe��'��@��V4�J�¶,�PH�RQ��Fܰ�-�9e�4��9'> Mw׽�kԽ�1P�'[�|VO����x�V�3�jr�ҝ��B�9�,�V��鈩Q��|&^�*deҢF$�7��A[����Yb��SOG�L��c7�2E�x"���)����O��3B���ĝƬ���W�!:����0/�������UK��=Qz�6\�4>��h��(3 ���B�W���:њ�2�c�3�ze	���ߩ��?X�����J��o-����Գ��p�T	 b�v��p����0W#������I1��oQB�����]"�xwp��a��x�X��J�l}=�1o�v�'"�/{�<�H��;,_ì1M��^Uk�b��'�? E��o��DH��,�Æ��m�
�<�TZ ����L�W� ��Y`o|-Obnp�V�����ڏ��B�lr�E�4\�-�>����'���W��]����|�Nh0H�~���u%�t5��P"�����+KO�l�H�ه>16��`��$��0"k�H�8; Nl%Y~��������\�pd�[s�rK��#RT��w��7�w�܇o7�ɻz?@*5�3A<ռ��g�M��ɕlY�b�����U�t'h�4���4�;p(�H��ȹ�(��q7y�<Z[������������1�U򛼣����^E�g�f�)gF��XM��/d������񐛳D�@�O�2��T,Vw�j��drx��MtSS=)"Tv�%&��U=�d���e�f?k�{��f�2�ǖ�	��bs��M��YJ�`�'#���qfh�F� K*(iKJpLwJi���t���{���,W~���cA�]�,�+0o���������[i��>��a�<��?��s���`˹T��@ip�3�Q;-r�sNj?*�����r��A���hy��{oX��
u�Xu:�TdtZ�0�w4�%�g�#x��ޢPrK�z
�zpx{#e*KI/�@���lx�S�f����X���ʬ��>���<���M�Ψg�y��!>Q�A�z��K�����3����>'��q:|E��#$]ի��&����c��^�|���6��R��ub��j�0����<���0��Pr��%D��?D[�"*xmzM�@�(�����bjh�`�B%7���9��۽od�֮/�?!���y�b�Ȉ�~ݦ�g�K�����$K�c0%�e�]��l��!���/�@s��X�$�#����G}>:�}*�i��s�{+)4�r�Ri��HSמ%2+�yW8�~q����ټ�M�XN�@��@�pyT+Z5�5���	9\C�C;D}J,��Щ�VG����#��qծ�%҆������P��3���Q��a�k�>�/���D*�M���
��O�O�rDS_[M�f����/	����v��s���ջ�Aس8�tЌeG�������Q��B����yk��M��T���j�^�O>Um}�ȵgC}�:u�{A�b6���i�oL�(0��&���^ ����z�V����5�ٯ�Ո�WgS�=��ʽ�"��3������t�ԴʷX���}��U_�x�	s�)�v�~��\���xy�:���!@�G�>����FB6m��Mq�?n�K�)��D9-��<�O?I(
�{Ν��4.�M4?���lR@Ց)l@��/si�0_��h�k"���7}�Z�d�|��p5�<�.��0�����P�����Kr/�c�N��'�H#��!+�TV��:h\���SaJW��)�&N������ԑ*t�5.�-���,.0�L?��%�f����Cnag*$H�����$����(�wEf����$َ�1 S|�UX��Ρl$����K��w|,|B%���(q�O�~Q��Z��7�6�/�sWs��G��~� Q�~�BP��s����Ofɛ}뻾� VH���B��0X�(젱N�kH��(�m�c�bQ��G��rR]�$[�
{9�;�|���/Uъ�����u2�������`̛��p����]q���Mx���G0���1������E�$n Q�����tn;�da*7�C�	�&�Tⱊ�f�I�6v��)����}M�AcWJ� ��4u/|(�1�y�x�J��S�m�F��KI�R���3�y>�i��+�v�5�Nm�@UZar����OpX*-E:5Jԇ�x��h��ݻ[+�#Ecl���C���̿��	 )�v����Et��g��\�!�˒��?�/�ĭ$���+�`B�/���,�܁E�s� W��0b[��#�� ?6|�j��x�7��k;\�%Fw��4RW�`0]��#�I�����Y^P+N��)w��Β.W�ũ�8�0H��3b���4'@:��?n�Z��X:�EM+�EP5�,�.���5�z���8�B��R��
������/g�8E�EnxpNPZ�����^��9�Ͻ�����	���(�{�܃��'rp���j{��v[���%�Hm�[�i�.M�%j�A_<����٧��/�,8k����]'E�'R�:N�i�8��T�3HpMC2���S�\s�<q���X��+��o>)�_d�x�7�j��|��]|�r,�Na����AWm�O\��ro�M뼍���ްDR�A��k���_7K\Q�\����R�wG2 �[�
z	6��׵g�xv4��Կǩ�朋,���Iԁ'�l2�@��3�S�2ud�� Z�-�渑�=m��rw+o�&�x��7�夥�%\�����6���O�`�J��t(�	@�C��am�o�Ya�2�m� B�:7exy�:�3e�z�œ�,,a�=�S��7�s('
w&pN�]�''r��@�A͸M���u>��I
�����m�&p�J��{�9��B<�.ۤn��Fv�h���S��B�ׯ�ߵp;�Y��2�ݣ�)�f�f2F���9D����r�d\ ��$[]:�|�����j'n�&pM����_��[iT�U��U1��z�	g����;�$}����n#��Y�IY?,X]E�^UJ�<o��):�Vγ�F>���먓 ������t��D/&�]����	鏆Z�l�t���Z�]�M�x]%�ǫb���dJ��C�ӛ�jS �Fo
��;�q��Cy�������DS��Z��U<c�PO�z�O_�v�|%��\���0Wi43/�Z�)���41����gGƕ�%]u��Ε���_��k���*��;Q�|#f��Xz�ư�ҊO�| �h��`�"H�M%S���6�^e��'�陣�T��{I�⍢�X��	���!^��)?Y���d��/���E����)jq=uIA��c�7V(#��[��!�Hyf!�xc�c�����~1�p��,s�9�v�u�B錍ݲ^���d��T�'0=q�#��B'eα�G�^�P�m���kR$.��jn(WE�����DX�iuq���`��!p-ߜ�a!G�!��>��J�/j�AFf�R͡���d��\�-D�ar(�^C���!�N<�n�Բj-b����� p\���E����+�|�w���;��8����݃d��l0�=�+�_�pɉ��[ɒRz[V�w�-(�� �"�MaIExN������P�c����ajI'�$o(��9��
-X?�4��	�����TGpz9$%��*G8�����c��ln��a�b̑�]/Q�j�?~��B�	�3��$�:Ɲ�&��>��EQG��{㘋�G�"��4�h����P�<E��6���F�)�<g.�&v4F�U�&�\���ز��ÝFŸ�3��)Q�Y�G�ȏqw��Ӻ��� y�Y�O^�Φ�����I�+�K��!C��Xќ]������n�<�f��F� #
�7��T�rca��_ٖ1��ނ�'��:�� ��Ig;�wC�1����f>�Zgfd�S�iy�����n3��o�˙h$���`�5�+�S�@s	d�e,Y��M�Ta�u*��y#/1dӭ��h��������Z���"A:���ֲy1M,�e�Wӱ�p��z����N�5��$�s]�GW��d��fg�/�LouM��9�8��#{K�{q����_#�cR@�А@�'<���G!ݷ\�&!�>�\��+q�����l��	[��~vCCK�b���ɻ�_�$ɋg�pYM M�j!]d��u`ks�P��ED�x�ǌ}xMmd۟�d��L�%�ԒYb����
.U+�K�����x�y�X�P;C�`�f� ��B�Ѣ�xm��H��]hp���ZǸ~��;_o��N)a�*�G�n
�N��fE�s��B�HYg���V��x�f��_�+r��
�>'f����f)����]�W"3�O�qőn�4T���Y����`Lz���xH������ݭk�~�=��2l�wA��yh�+J�T�
� �]�D%�{�MG�9��.��IV��̌ M�K��<��%��ބh����>,�g��%\ K��(��	�۱���,BE��������)P����9S���e��	�RԄ}穝U�O�M��c��%p��m��=��M<��U���~#�W�L���Y�w�fL�N89d�T�/[H��@��R�wo��&g���'{�c����Ϻ�t�g���I��a�+d�-;��\rj8X��6��)�9��z�^<ӡ
z��~�B�Ӏ�+����׈2	���P;�7\���]�N���B�?���H(y�c��֝�W�)�����c;�<h+��1�y��Ɏ[�#�QJ#�P���&�ґq��]=7,B����k��HG!K���~�o�z��`<͚D����>\��������/��d���ǿV���A�Sz��Þ�W��ʚ�D(�f���B �]F�i$6h+Hi��Z/T'M{����`$�it	j��e�K)��P�˜��n���]��7��?28�5�wo�v $]� �#�y�O�&"r�:b��6���tb�~����#&ڡ�J#�Ԕ@��[�uxԏ�B`'����VL���pذ/�m?�o���EZ�?9�a��,3Eym�`Q`5pġEҫ2h˂�A^�Ķي\PmR!����ȟ��KL��V�b�}�>z�B�Ǔ�e��:�T��@��VE�E��/�����m� �M����
��$�)���s�GA�/ȴ!y���R.u�6� 2q��D�ZY$,5Id���,��D�a����$�6�}?� ��v���i��vkD&����r��	�`�,�$���ﶵ������UQ6s��2g����r�}�2�]����F��>Ljx9�y�g��� �����\�P��&���x;�	�%�G��gv�Z�-�{r�G
;���[��ń�i0�w�Yi���3+�"����Zީ ̅�/='F�b�ICRI��]�)��G�3�]\C�:m$�������A��^����x! j9`;rE�S�$�� �{0�}����)j�x��Ę��7U'"��T)iA�2�Y@n�m������{�%�v��l�7�yݏ��>Lb��X*���va�f�����d��y��Dd�("��Q'R=	`I�r��pQ#X_����+>�_�x��͎�\wz?*{>~�͙^s1"q���2M=a���b�m3:?^�$I"U �<֟q�bŪ�����/�G��$"��*.��De��3��p�b��F6�6���⌕0g=w��#�6dܕA\��8pP}52isÛ{��9G��>�"��~�84b���e%>�W�1YS�"MA� �l���N7ș���5'���G�G6��.bm���V�3��l�'�c���� ;�۳���� �W�CV��b���!=���γL���f�TMҀ��O }��x?�0�=��V�C4�F�
�1�f��2�~� ^���	��5O_�vI���7�4��Je�[X����g	�0�'����B.'����j��{�Rd��9&K8'�R����Qٚ���2��ۈ��x��S��iϥ�@'�Ø�]ӑ�,���@��3a	��*���A��5�_}Ԛ�u=��M� ��ti9ҕO��!�6�}?M���^��C�sr8`n��q�A�r��bP�������޴��� *gG�;���HE����ձxT��A��-+].��G���J���:}�`9��$�_��(݆u#
<+Yv���a�Y��&�e�#�ԞWN˒�C��Bd��xF�o�u]a,�Nۃ������(�E�Ia^�EӀ�?/H���ٮ��Z0zD��oJ�?���/��cL���A�t��v�c�˦��c�?�֣��8�p ;�/�������}��x�=���	ݽbe��K�HTu�m���U$�k>uu=�[7���2�� �����)@��4N�)�W1��H������ +�^����7�?�k N�l�Z�{��w���bR�2c�T�r�b�F�"�ص7�$�z��j����'R�f���Щ�a~�����O�b9�w��B�`ub~F��jPMF� �c�7�J=�x �IK�d�[x ��}y1�!9��T2�bu��%��@�#�ϓK#C�Gy���A��҈���ԶXS11Q|��3�l�ZV�qTy���yv)�. �M�>�$O�)0��ZN-��_����S�LMc_>���q�X���g����{{͓9������	�M�s4��7����ѺI�>�V��@}L�'f���\}~E�W*wIŤ_���WT�`0)n�	���tC�Ś�`�޲e]�b�2[աo�%A�yG5,���zBY���{LYr���&�vGݷJ���q���s�"wq��"g�ؿ�P%6ڬ.�48�Z�^&�d'�ͧ�0����G:YơJ�@��u�������_�.$ �ɍzh���zd��G�YDe�e�ʿh&�j�Jh�8��e ���(&�}Lj��W����ֲ��*(Fؕ��+:X0J
�] ���n�M�s_R}CϢ�yʐ}'��4�,G���rZ�r/m�m�~�(SR��X�߆C�B�	�q��|�'��78�S\��fw�Pɔ�X�40�����/����t¼�'���e+���,����ؾ��ݹO)&}#����Ocq�5mRW�7�*���"C<^C��?ti�ͱ~F��`�ߗT6��Fp����w��R�F�G�|�.���{@�2��K��G�%#j��%�F�/H�bǤg�3h���ݰw<���	�~��/�%s�9��͊����ώX��z���҉ö����_@��E=��g��w�L�3��,��h�Q$�W�i�����X�p��p�k�X��,�ק1R��S?E��̻,"��#�{��Qz���I��6W���=ʺ�v@[�H~T'R�I3{��H�g|z�|���T�3N�ۖ"�,���[A�6��[M}�G��z.���S%����q��	�4y�_X{��}���D�}�&/D��t�|�O:���T�w[��@�%��G�����B�_��@��0)xr�I#��Ea>�1���#��1(�t� ľ�/���\W���6mN3��3|�`F�Ԁ�5��u��^O��[x@2t;>XJ���L�-ǔ�c�����,d�[dVp_'Ç��J����L�D��_�G�n�g
H�K�j��)���GN/J���P�Z~�>��g�8(��7_FQY.��?e�)��#��7�m}�*�y[���}l>���ʗ�����j�%0����!��e<d���K��
���%v:~����ƴ�3�Y`� �8�Y�,����l0�L���y�v�fü�n�?Z�q��.#-i��2!z ;F�J�	W�cT��#ಝ<��z^�6`���p�hU��<9��1��E�#��"�
���c�2C�]WԷ�� ���"�K�ĉ�eZOD���xNC��z���Jɦ5�bq�UZ�����/lO%�y\�v���P	Ĥ�s�����U�o�v,�S2�gG��:㗢^��o��~�U�'.ȑ������J�^����{��Hξ.	�{�L��i/��Z�%���3tC�':��7+9@���'��d���nQ>�9@D�H�X��Af�+�����J�����z�b"l��<J#��Ct;�;2��N�@���[�s?c�[�]��0�k}�,Z
L����ȅκ�� 8;�+Tu��+�~��q�Oo� ����%�6p+�/%q�9�;��H��������� �I��ş2+4Macw0>!\���]��1h�h�s�o�G-��o�+w.�8�\�c�x�9)��z'\�t����r�wS�-v��S���R3Û��6�#E��nn&�;s�Bu�X�����Qx���	^Ԑ�V�4��꾯�n! ��VL�[��~9gW������Z)6�_�.%��)W��6����z��L�w7Н�JD	��V����3$L	p�NƩs'�	�s�5��>>��W
��m��_l��z�S~ 8En�+ߎǆ�XO�Ef���g`�����'�v��AZ��p�sV�ÝUl4f���Wo�>c�dY��ڠ0s_ʪ��"�ya�V���	ÊD�3`�UU���B��n�B[`]�FB" ��4��7�9͌�x�5�
�VL|9de��[��p��-�E������w�m���.�8rTo��&�[.�9�a3y
A)B4�����Ԋ�7<g��#$���Q({�K
Y�m��(R��"��焪��,���&yb,p�:��_���ya��:I/�������<��&���8B��|ᘡ��F�_�j�1�^�E`uH�hz郞u7�1_ě;����d-����u3�� N�r�̫����^�	ՅR��ڑN������We�J��kN��6�1�+��͈���g���B���;�Z���a+;Eȓ��&C����~�7�X����]����C�mV|�%(Q�ҿ�npaːm���`7okUG�d&,�Ǎ��K[���� �&�P���б�;sL�i1���Qȣ�$1�	�Z�+����(�ږ��<�]� ��8�7����@�?A|�Ve��۝�g��ԇs:��{��"�uE!�:Dځ��N��z�	�/i ��KZ�9�H�Q?갯�����j�d0�/+�KM�UY͋v�\��� չН�t"��YO!6�u�z�jc�Yo�vp�ԭ_������ѳ�K���U9���[l�MZ�y$��ģ������>�|��Km�������ߏʭX<�@)�����M\>���Њ�G}�����XKӪ��J�����T���Y�9��Fd0:�Ȱ)����"	��\;G�ɟ=���1ɏH)Ouq�Y�2
U���7���-�S	�pB����L؝����{�O;FI��7�4�i0ۋ�w�Xqb���{;�A4��(Z}�+�Y[��e�^C���e�nT�u�8bE�ď�����w|�$P|I��M&>�G:}����W�;-�@�`(~<��Py��өW��z @\4j�_�{�n@�8yy[�"$(��+Oc���O�'���M��n%**S�����,D{��s��j��X���IEL��o��q%;������{Z�
���*��׏��R [P0|����	�"��S�"����O�<�s䕯�.�ʤ�����e�DGen�S��O4�����b�@a�j	���:�r���F��EK���x>U\�" ���q��z�$�sV���i�g-��!@�A_�L+I6��wO���>��{	�
iʥU~}�3n�S�~�(���{��y�`/�T~�8��qq:d����Ԛ��b�뷮#���BQ�F�~�(ٸ�r��}���Q[M>U ��5v�UP���{��f�����.�oV��P����C)�~�a6�����lހ��{�##v�:o�^i�'��ΖxF���\(8`���F2)c4�ߞk���,f�����}�VN�O@�h����
:F/�p1#�̟�����iPp3����R99"�$g+b���jdPY�E�8�r���:?T��٨F�������V/�ȍ�#�Jw �U���V��A4�a�͍W����H	Vc���Y���h��R�m�1����!�Ӕ0��S��m7_��i俀a�&0bs�c<з�V&��L�?��Kg̀��`�Yd��-M�?��J�˵+E7Rw.� � ��Q�3�Մo�,PW<قU8�?f��WU'مS�PN�)s��i��ca���[��1����e��E�'�cSZ�^7�v���ٱ�:?�/K��߼�Q�B�L3�(@%��	U�~�O��Q�q��w��[ъz$�Q�Ӱ2+C��P�� �>*� �5���>�7� �X�`���o��05�eX�k�6�-B�`i�pT��gc��^���(ĊN#�A�!�h�1:	�t�υf~�J:&���65+�q��S���1��J�ΕhƏܥ���)�"�L]@[�ӊ #p�h'�c���l!Q���.�&��]�+k�x���H�܈��y�%��+��H��p��jß� %N��2��.(=A�B�D�x���?�#ƙ���\�E�Ůh���e�� [&z�9.����5�YW'^G �Ӥ���v�ԩ��|��h)����OO��u��9�*�Q��iW�r<{^)�����%��!/�4��"-���àTq�w��q���W��ޑx�k{��;����H�A�2p�V7�ވ�6fIV�g�Ǘj �th�soV�@��z8d"�b_���=Ⱥ�o/�]S���Q�v$�V�t�����+�v?s6�2A&�{P�;��-_����7�����Ʃ=�`b&�2xS��Z�_�N�L\L3��}�\�d;���??FH��+l^I���Ie�����z�-!8�i�W��d49����L��߇z�ɠ𑻥��$�����/�%F�z�><����z��||��03��7/6%��:��&�|�Fl>�=��w�����iv+b��h��#�t���yZ7'W��;Z�Bi=	���o���˔M��0��L-,�iR�%��f� *���J������?�@v�xǹ�D-ٸC8�}_+_[��s���	i��?5�����������}�J�B�ؓt8��rs�ۊ΅k^6�4W/�Ꮀ��g�qAZ�����b`�.�C�/�U>6������x&� �Q�)Ȟ�~�}�d����;b*���ɳ�����ݘ�dY30��L�"�V<<]��Ŭ��,�mhH�&�t���~��Is 2��a�k�ɔ�w��w���1�SQ��yQ�sO�;�r2����+i|0��f*�,3/j(daz�qz>W�V����0{N��+j���S��%�����ʁ��,�<W�W�2y����,`c)�Ⱥ{�uzm�c�(����l�FU��\a �Ʀ�g��û��GE6�Eʫ���X`�������W6��գ�,��ۥ���r�|$!����hc�A�q>��>Ws�֯d��WB1��8��O'���� �(�,6ێ�(�O�[�0P�� ��Ac���I�G���b��ji�^XI�,�g��=�Sٽ
�Ȃ�-_�"[�*���Xq\m/2;�H�o}mm�n
��f�)���N�[�]\=����D�ɨI��q�ʬ�j�y�`^X�����e�_���Yd�x~�azx]�Į���ok̋=N�TA)k0��� '~���+�έ�%n<&K��`�0n	������)YN��ø�f��h�oQ�G��C�'EC�Ag����l7~0)���V�r�KJE�Wm���Ԁ�:�S�=/�{/A��QU��Z��= �`�� l���gX�n'fE�Q�r���%[ڃP6�����+�bWp�W)&J�E�Q=I��
}Bi��]��rN�C-M3w��ه"��
D.D� F���(�O��ev 16UH��q2ZCd�hK���h3t��ބ��0���Mg��F�a9?�+���i7~�D��!��g9
~��%�/�4X�S�X��5DS+����S�ANx7%P#{V�U�Qӝʮl,1������ɪie��Ѣ� �=V*YrݚK�����X1I���E��z����� I�lL
�9S|գ���=���sr?�r�沽'�C;�3&gT��2C���H,L���*����p���
�p݇sԚ[}�8[0��#�pw�^�^Jh�1�ņ�Ferv ����m�eG5��G۹��P�~�峜O��6E��z�l�J�D\C۬x1�f(��ݜuL��3�)[���J����"���}��*V{Ǟ 	�&�[��0�����{e��!���XQ�V�kw���	�y1��K�4��;��!/��rv@@\����j�ݯ.�N6[�r��ԞطVn$�n�n3�4biV��b�4�h�9���
!�@���
���grō��7��VXe�YE>щ�뺇۴�`��Z�If�Id���j7��9������
�J?�(�`l���ڷ
��퇣iJS/ӥ��LuE�&�<-�^�˚����<;�=��1�U���t�����:�L8�{���>)7�&�lM�:�7Kd����eծ��YV��O���t��� �sk�=���"~���\�z�����K��U?g*��D>�˚�)2�@(�D�^o�{�b������`۰ͥ�����/U$G�^�S� �ju���ܼ�k���PC��)D�?w*�؈>g{�)%�����FK�ᲂh���ũf�$ߛG�6aN%�9hyY�sS�R��`�1�]���9/A�!�[���N^�e��؜k����(�jP��S�"r�K��L#A;	�� ��ǎ��H��?��'RR퓓j�(���4���ׅ{&dO���c5v@n�L4��^��ؕT�
<�',?a����|��������Nb �nꓝkUw���(���A҆ܛP�P�n��s7kP���c��BB�"���ђi/j<�8A|�y:�g�s�W���}�y��f�l�N�䚨]��y[�ui!��L>���*�,lwK�5���p��M����㸔T�l��V(�~��Z�u���ŏ>0�,���8-t�񀧚 `2N	�ۉ�[Ti5#�I���l���qN%�P �aT�$`��Rɓ T��j��xP���00���z�r㭛�3
�����	�/M��Oq��s�����A��M�Z�-0!2�UğnY5��� lW3�X�T�Ա���3~�����?���p���! VRC�U�I���Ņ���w��E��ٓ��CN���u@�b��_����m�H#��T8!���7�}�F�������&�jg�zP5yѤ=ax`կ��4�2O2��MM��u��֐�u�Jӡ�p',�u��N#LO�]�~^d`���{4�*�ߤռ!���e���?��M�B#J���)?D��l��4.l�#s(����}(�B�����^�h��B�ߧ<�U"gyVO7H�*}	�S�F�Z���q��D��͹���rt#�Pc�\�cd%hlc|��E��fO��|Z��;NBٴ��Ķ�_��2�^�Sa�1������j2�Kè$�0��Wy~��Ň���#��o�v't���9{��'&
��*�ҐjO���d�`�W�L�%�B_ux|R�\������L&�V���{W)�X�C� F3��\�x\?��v�b�[-�=,&��a��I��M��SX�y,�i�]���eK�c� ��I��M�<\4�uwM���s�H��'�~�|Lw-�8-��c9F����F�K�m�OoX�U�.]UCQ�S)<��7Zܾ*Ȯ��G�����2?��Eer�nȷ�W����L`�6AΨ��`,�b""�Q��!�.[D�*��$U-����rGi����>1(6�7��{���h�E�N�}$s�e~���鄋�=-�j?ze�dMA����<��K�Yh
��'⯈���㡁�P_�q����y��Uv{��a%����`�}�{�k`\/��D�Ƶ�M�`:��xV�d�P�B~��e��7��yy�Ò�T1PT���į�4x�q�7f=����l���I;D�ߢc�Bi"?���X�2�
"�I竰�s@� �� ��뫾03Ð��hH��' [�:�~<�>�͑��q�8ax�>��ZB(���W����k�k�O�wޥX:�c���}#�	��6��d�䙹��w�?�<<�=�iD�/M�/X���L����k�pXw?�r���!���q��^*�[ϲ�@o�_���
��ib�1�����N�Bہ+�qɑ�.�����j��Ѱ�+۷�y���1���]K;��m_`Wn��(=t����'�����d��YD�^Ϙ/s$'S�5L��&f�w`����`�VP����y�{~����sX�sk+�v5��2�� 5 �V_��F'S�/�1�U���2ꭆ�oZű������~.�Ȝ�'��	����̫I����1O���j&-+:9��t��^�r�N��+��fx&��O8v���kUcg/��+��	υ끛��-�[��o/�~�5Kޮy�5d/ح0ςl)7�T�Q�X���N��ܲ��DHfz�^3���|�v姬�&�+�^��-�<Ό�G8��fq+&~��e�xa�L�զ�B��eyv!-/�[��/ķQ<�pw�X�[�)vO{������'Q�K���#���St��H"M�	��Ȁ�*��1נ�7�S�@�w�{x�Y���Z�^��{d^N�����e���1���w*p5b4�q�������w�����Ϝ���2��nb?4�#R��)
�齌g�`x/���-z�2�R�p@{4v�Q����V�������W���dͰ-��	F���gaC��b�S�5��&ӕ�i2��9�����z�c�a �)��U����6H����.�y[j�H�qQ7�9*QC߭��9�%���o��2�M���Jո[U����{�×�:D����Y�٬H��9��%Ђ��^��Qu�aP����؁y�.�s��n<����9c��x��A6N|󡧟���i���ԝ(�g�|���m@o������D�1Õ�r8? %`J��
0��,�#:��ԯ�T2+�Jj���IQ�.�lqV���ru�������b�)�ƈ�zp�!�|�v�{l,x��ж
�M`$�}��+�o
���K�ДKƴy�~���$#n��Y+<2����d�;4�B$��s���Fcl�uo�'b�����E�
�͂�A@(�|���=�p�=,��3���!sy�[�?���U��{�{���툪Z0�x������a���W�m�a�j\�swP��hf�&4U��6�<���f�':�������+n�O�t����O�"�↫I,��C��FH��*����u�@ͺ��50J�Ŭy3��.R\�t�R�5K��r�u~�ށ�L��8u���E����48j�u������W��Z����<���6{�.��ԵU��ZIb1���.a$X!z��D�3�j�`�v�'�+��5InHt9P���SO�s]h葡ɔ@���8�_w�G�s	2Y�~a�7�ۙ?͢��2I�)0��K�k%�:�h;88�}:���'�Yr
�,�y����Q����A�U2�E�ڀI��+��$ik|��e��Κm&l-����$_�4v�\�% �|$����/8�'?�Ĕ?�V,:i�O��I���:<5�{A%�F�@_���c=D��^�f�r�$	�GE�Cw��Jkk�WW)��!Eٙ^�.���cN���a�M&v�-S|���em�;��n����Oƣ��Z��ą�z�.��a�%y��	�yW(�-��^ϣ,�M	d#-���/����P�������o�[me=�o�h��`�_5{AT�nMsf�p��v/�s��������Z����Q8�A�@�|�����h�p~[�j[�s���
�<�����^�:���c��݄�P�׆J��3���Ľ3<o��0K�і�E0���\��8�;�ҏ'.�2��j�aǓ��*j Y�3�{ѓ���WbR���ʊ/�P��OVf��$}~���p�K��`�!�Y�i¿���=D�)z�>�3".-��IM5��v�?wk�Sy��a.�������7�1�F��#B����3������C2�p2�Ƙ�f��9;�p!�یXrgW�"�g�P�b���C8�H
���������W.���cW��[����n�	Ӹ�a+��~CWT�nU �m0�V��\������Lݗ�l�\��*¿��X1F@ޭ�d���̐���T�o������HJ�e�����3�D\���e 0�E�5[��T���j?p�<��(�Al�]Bu�|�c��vu^�\7:U�%a�=��Yq]�_�q=N�N�H�ľ�J����2�%z��=[���F=��wC�G�s��G���ʆz������'���b̓��+�s�8�Mk�l�f2���Z.K2��x�5�KM�R�	�<����9yGTm��;o�5��p�=?B�-���Y@�G?���H������q��QaE�9[�:�C?���2����O�����_�6��7���w�`[�-M
��nd���y�*a&�!�}w1+x�%�����JG�ڱ����qS8�^����(N�)j,�{��o�6Ӳ+8'� ����ۻ�m��#� ������	�)�S�+_;ƃ2�^¤p�!;B�Aه��e�XY�M�Bg$���򤯒�ԃ���=�#Z�=����Jr���g��m=�l�&躤�jG�X��x�������Ю콚����~�$<�6�wd����O$A
�k��4�%�Q�����#2������V/��OSײ_Sd�Ƚ'R�����M��v*��Z�5Ucxjz큅~.����ĮbՏt�A��PT
�[�d��(`�Z��7!��n�#�c;'w���$!�G.�=l���\�~��k�z`�� ����J]o0���[T�$�H k��o���撚���ɻ��So��{�-�F��_Z��R�n����8�%I�����0G����T�T�;�5�3lz��Q�����%�E���'3�Ա�ޭS�t�c�@���l����8��c��N��!&��=R==����y��Z~B�}�]E�X=h1DF2���M��{���!( ַ��B��Ԍi�8�#�)�'��!qe�^�х��"�%����,���8dpE�A�nl�9�� Y
����@��2��WZ�	�&�	D����1�Kl��{�|v��U�J<�F����|��C���Zw�^<��z[IHC� ن�	;쇄�P�RX�r,֨��+=F\�d��J0�a���Q��{�!2/&qL���%��Fv�������{�a�E��v\>�0m�|����l�ۓnHpQ��:�]O��u,^<�ZLʞÂo��Y�k0��-S���Dk
��ɨ��l���Z*�F�*�ݮ���u�}��q'�Sr�.��d�sI�M"���ٍ����P�ɛs,/��a�y(E8���JT26b�F��GW	z��!Wg��thv�<A��8�n�C�a5bX^f�i�(����ǧ��7����(�����r���ӎ�d�<I�_�����x$ߖ��tnV��bs��ue����-\��z�u{>�W�PHZׯ��O�'��E�狸����'\�7��ɟ2���I���){Ƒ�q/����4D�\�r֮5�H��s��_�����6�S��:DT^��Re҆�y
b�'߄e�|t(����词7��z�5�$��56c���8��R���p�s��/a�}�s�z�h��a_�Kw������)�d�/H�w*geP�@�'��T��p��G�Widf�&Rq&������� ����D�=TN�$C�2��'$+�<���Ա����aSt�+�����7��\�L|�o�m)i�x��:�I��!��\+� �E��c�4���8�4��\k��SP�+&�n.c�zn�;�
��~��7��䄎'WK����昣^uv+����S4�f�d����/]y{:�"��Xoh��cjv#B��I6(#W����!P�r�H ���x�{��uA��\{���N��Y��$LϱܵF(��c'$�גv���u����.8�G��p]�z�|��Eh�XKI,eF+�h4��ֻ������]03Ë
�K��
�L��`����@u�C_�^C#)��P\�9��:cG���u)�&�[/ِ�Dp��v,����-NS��Z"k0���1
�9�R�s��tG�ᙇS�~�n���3NU�}e܁<�i���y��oG� �����1c筓l��5�b�j�A��Jf��ρl��Px�7�0��M��`��I2�Ƿ*i���sJ�#/���J�+�7��8��	TM �+�����~b��	]*9�}g�?z�����4(�ς�9���"��{��h���j+���������8`Gt�"�@վ��4{8�++C0�#��qh`�0P�e h c��ir-L:�x�ŘՓ�Ϊ�]�g�M��Y(*�Fw����.�z���d��T�����\������p�ꎺ	=2g;v��=���2N�� s�����6�kt���;E*pf���Bt��nH]?�1Jo�q�����6Ӗ��X��R{�*wٜ�S�ҷ�ѐʻ���ČC|��� I&��U��Bq	7� \Ω y �S��X%�X�6�Kg=��г.��먂�����,a��5�?�9�B���个�r����φQ=�9f����
��B��1kW�jV/f�]�HR�,F�T��}?�_?q�?�a?���8���܄��73�$�M�?r՜��q�d�%����_0C񡷓���inm�v��v�
|��
p�����lM��!�����ޯ� ��)��؈(;��]�"rߴ��3���G	��0:�����+QqE�����!��D��#;���R�0���
�c	{#&�t2o��>�M���e��~*�@s�x�qm��7�HZj�]_�/� ZL�^������(����tP6�YGꅶZMw�=��4<H�!���D�E�ʱZr���׎)0@�B����ѐA���*��Qj�N�P�o{�_�;y'�*�W����`���a�*,���$ۿz�����;�N��YGc�\�
} �`��+a<�.Z�!O������7G$�'tPr�:��r eK)P<�/�G���՟fB��{�,!~���ΫR^��dC�kH�f*��h�_���i��Q2gcJ�� O���~~�΀od:1�p��Q&�?n�uWuf��8ڧ�U���a J�$��&�p�"Be��p��'��KH�$�F��<�9(���]M� ��/}�'��I��R�%����N��{�\�>f3�{ÁRUW��4M�~�=�"'�,�כ����g���):�����z֡�Cʓ���u���xq�Qa��o4�������歷� ���I�1%��kN��B�oD�=�V����<?�?N�700[���}���7���d�*<���D sm8�o�}�bmqp5=���D-��ٷ̷�Y�1s����|)"8b�9@�����~đ`jb����P���mB<�g:�������"Y��ڷy�SC����3��S�M=7_|M�_��T� {�X"����nFU͞:���Y�/�f@�ր�ķ�N7�� ��p5��o�Jv�0�I���ˠU�A{"%�iz�)�>�I�{���W]ي�m���$D��l�֘$��{��9���|.���S~陚0%�N�ke���N�I�Ң?b�ϨӲ^��ІdA��r�Yw���熂֐�3�Y|+�e��؉�^]8����A�-���_����~���U�w��Ķ�)��鈥WW��8� MZ]�r�0$�m*:��(Xu#��icZ^���.{�}k��ॄ���
H��v͸���01Q�1��OV]*\�~��[y����rVl�FI�Z��-���r�(�[�o�d�����u�=�إ��5�E(�,P��Epm��Wl���<@ �g��a<��������K��X{+���D~6�
�릯_7�{v'e8�� �]-�lXs�cG����Z�=���]�u^MvsA��}��eG���2��"��c@��v���W�x���_��i͟�	�
�>�"�h~I�0�DG����F$9���B3(� �۝�~�&y #j��1���:q����K�(�e�Ԉ��#A~�%"֜�V|ٵ�(r0G�c�g1-6��rrv4/���M�TW��C�{s(�VT~n�ƛ$&_���*f�&��-9te��h_�?šw�г����_̟�m�<�G�;#������bƳp옧s6,���T��! �z��Wz��� ������fC9%E)N�tF��a[�����^�H�$�S�$1��{\,L���p��76H����ë�&�45��+�Z���L��'��{-�@��Y���ȑ�Jގ�\��'P����k��a}0����]z��se@!����d:2���i��v��zQ^�3rk�ԛK9�RK�_^����x{�J?U��:��f���sȔxJS`܇�(��E�ĺy4E��*�q$���澁��z�;(h�t'E+�6xh�ʭ�b^kl"g(G�0��}EJ�PJ��$^i\��%��=�_��	,.az4$v��u8�Œe7`d%H�H��ﯠ��D2�ۚl��}�IEo|6O�:��+��^12� ��Q�C�N��Dn^ӽ.[i��e��(C���8JM��oŐ� b-|��y���1AA�~'i�P�{�v8�Cҧ0a֯�s:���9J���W�-�+��sL��=���he1qm�q�J��"S�D�'�;�b�;�S�.�&p�2�}Hly�y����A�&̱8���Pm[�Y m6������5h��8��{O��a�SB+T��X���UHΓ:�g�1��� ��m d ��.2p�`���#��Lc\����� HyLD�䉜�p��)+K��n�#�'��Q$��D;���b}�Ǉ�n7�v��a��fU��] ���9|$�<g�0����}��m�l�:�$�k\m���t�J3���讔V<��g,)K!�y3Q\V�E[�n_f�TҶ�|I�l�E��oĢ�{�ݖR'��iP/�'	TQ���x�B:�a��{�����A|G�{��Р�+��ez��5B������w�)�ii�YnQ��0qf)|O}���%�mػ>�Y��pVHm�K{�#�GOU_ž|V�t>�żw[O�	����ك�mO|��ݓ#Ɛʭ2�N�I{j���N!H->�tGh���į�L ��fs}@9f3ə��T��䍉��d�ĺt�ॶ����c�fE8MWի��_���~cI0!y�Y ��w����g�i��Y�_��e��($�oΚ��o�Ba�l�E>��v��Y��I �.r�W�/O8#��ذ�>3N��?�i����q�8QE"�v�)Z�9����Y��Ke�㿝���#�e'q��5��&�#�(�f~E�@��&yQ�U�G"M�9��|��B��`=�KE�1Y�	���Ϸ(�:1 ��0�2l�Y��*�LBt[K�qvAߩÜe�������*HY�y�L�R��V�M���%]ܼ��;�G_j��{f���{
�M�:`IU4-��BAx3��D�z���P�ZG	�X�� Ӝ�/�4��X��8�����=2%e�&��8���k��ci�]6��a�3�:]tMGa*L�\���?S��B�h���6	5똭�XU��n��{H���4P �կ����#<�Jq�V/�+�&ڒ��9	%�XBٳ�;ҋ��j��q�D���X���WkPc�w̏�3��j
�SVw�Ա����R��*P������ҿ��qƓR��Z�H`�Q������)|�3C�$���,���+���%��3�_=��u��?y��)������M�F�/Y�y���$�L��4f�vsZ�p �����RX�r��m�}c�~�Nd��^��1���Ot2�m
6h+��gMQ������k� k8orq���#̀���'<*¶W����x�8���]�"C�V ~�Blk�Ґ�n�3a��T>���.�.3H �bc���GJ���(B��ڎ�"~�t�`Wڽ���(A%�Ѥ��Ȗ���j1U���e���_i����b����X�����*�R���I�!-6y�,d2}OW�} _�gt֖��~���a�f0�e���N�N`vD�h؁ܙq>m��@��$�<%W4n�˒�qI�-Et�ʛ#TI>\�OL�˒*-�הu�׼U'cI���5��a��=|������ֶ%ӓ��Ib��q(*K�f#�j��EJ|���W�ٿ�@L��j�r<P%���Z��P��Yϋd9���G]��*U.�X���yV���]�SV!������.���;�eq�����t̺84��X��yy��'���u�-�Q��͔-�q31b4��sB���'�lpl�
mR�mBs]�^7 [�O�FV���<HHr�6����8���ch9қ1cN!:?p5���B�j����ą�&s��&�?	�NF����B�O�e��W�to��ӐR��M2<6�krw�l�_����[��!���|�)���&J�ZW� �qg�)��=p�H�p/ ��M��F��p�8�O0}�_�a|7]_���%��vT5>��L�`:q�����3�*jr~���#���b1mi��f��@Ԫ���È}��-� ҿ; �]���w[�	MD��D��{V���k_R��W��r?��e:�++����VYS���9�lH��`Y�/����?4�՗�����m�~a��p��?yI�=�D�nYG���mZ��e���p����c�"�^\���=�͐˻K� f%ZS�yc������u����M������)��N���л����-��l������Wa3� !>���o�>6f�6ӎ����m�T��
����7}��=��b���P�
�5��B���ͨ��1g�p�5��5;����ɥO��Ӷ4��j�G�'��ߖ�ټMoVN�}��&l:~�qͦ�\�UႲ���p騄��U=�D��
��c�MN�ĕh^�M�Uk+���Z��iY���,Ǆ���ӿ��R^#�F-{|�u���d����<��J��|�B1%�u�Lǜ��)����GֻV��x��3Eި���$�i�^g �Z��B��Y��BIm���ǃ�5��H�eZ�V��3�y�N����tdV�cZH����;����������]y��G�p�)q1-�Z���J?C+9=�]��M�Doj��%�˲ڇN�� !YR`���rL�������]�,��%z��r���W�\����V�g:�����Zʝ	��I��������?z����u�o ���L:� Ď�`�T b4��Բ}՚jH��� y��71�4[��ˊVD(�/P�t̐$������y.�^�/�~o5
����=�ނ��ü��N��Ϛ>�WYu��6���涴hagT8�s�݅�� ��� E��q3�;��@�d!2(OQ�ǵ�5�%j ��nH�0��p
����_ⶅ� �p��d#Q�b'u��>��.p{�J�)���Seٍ7�՚��X��P_�w��Ŕ��v �@U�Y!s�^�ᬅ�&0��c%ZN>p�q��d,�	iB���'���3���B��!��5԰��-��1��3��e$<t���b��ۓ}���>�8�ruŊ�1e@Q��H�j�~C�/�	���/���aL>���o1J���_��{�
��Z]LO���$ �{A�~o�-�9��,Ŧ�x�hZ�KWS����ZE�a㽛/��5��M�{�Qv��w�����P�Գ���/���E��V<����:kq��J'����G	�ȴ�壽W^!K�D-��}%Ƣ~��S��]��U�c=)W.�|�N�����ժ9��X��ߚ�r�s��a�o�;@�fbb�\ܲSPu���wٗ;`j�tx���D��K��	�H�.s��o3�Z�j���	�;�Ov�ڪ��}ɬ}.�k��JeꆙƧ
ԼI���H6k/�!8�007���Ql=�AVG������C��s�Ŷd�W�ҟ��v��N�HH��@���w�^��>�y�i�Z�/L��Ϗ�؄�J��%�^{U��Xsz�O���}�M�[��֜�_��n:�o��O��ܕ�ՔAd������݀zKD>�y7��"]1�����A��u��W���@����"#�(vbQB�*���6sRs\|����X;�Ђ�8�q����xn��I1�Ez"�0�[�g��檙y�â�m�{��&�[ޭ戦{U�.�p��ܒ�F���2[Z�����gy�/�r;J���*��Vef�W#+s���z�AT�|�����&kXV�RCĶ&A�^vW_���z&��>8�敥�U~�����G`X��%�IP���Uz������ov�U�?��[î�ʮLw U��h�dW*Z��)j!�Ii5~R:��N�|i�xB�};ΉVc���ѧ�\j*��A`�${c��1�N��y��-Еx X݌��=��L<���Wҿ>���G��[�B��w��w���C
��\h�*�4qm�F���	�Ǫ6�2�4_Aa����5��I%E���<u����>�i��]�[�M�n����א�5�F��ߎ�Y�,G!}d��Wg?��R��}8m�O�v� ͵��]*a!R���fX\?����#�/�@x��a_X7���߃ȝg��K�_�qW�Y_��VH!� 4hIy�6��N\)0�<�6���_Ra�(ƽHAp�5��SZ�c�>��C����G�-d��_+�Ƴ@���R�:6�+�&������<�a�7��i��#4v\����aN�'��$`���z�{�c� S0b�ٯ���o�PRc�y��vء. Tw��!�c�l�e�l�9\*�6��9���ix��E:��~�W1��wW�m��`��flH��2�&?r�����1n�\����(�oTcc�|A�t�7�ɠy����mq��9�s���/ZA�\64�_��s�W���bl���F�;��%آ�kPc{Q��$��h`�p����H��uI`��S	߰� 2��J\	��<�$��5�O����]���	���M�r,֎���[A���SaU5ؓ{�5�H�M�֒ķ�j�Ֆ8��rpN��aq�;�p"a(���<3�W
�
������x�sǵ�ػ*����6^�>u(��rS�IGYR�I>�sZ)}X����d������5�h�գv�I��K�Q���]�D�3p �k2�AQ�,d��}��Ĺ�!��a��BK��V/��
g�7'�4�z:5Ϛ�yٝ�;�_���m�NP�6&q&���ьJ _�����8$��/R����52�yp�����y�k��R���N�Z������P��~#4��=���`��?`��yI�0�#oQ6�"m�b'<�.�"O��Q@=N������%��~�.�/@�@an���"�å�
�gf�B����z���C�\c���k�Ghse�D��'j�Y�����;�8�@�5uH'�4�������Eʰ��dG+�B4��O�N����&(�'��V�~HGiq: �'�{�Pp!ܽxGD	0��N�!��X�t��#¹���g��0vZ%��[�����C���1񾼒ر���X�-��x�F/����R��� ��"��e��CLӄ<p�d�2��/m�����MK��Q����
����M�5I���D�o�m���m��.�/��Qvat[��Qڇ�
jX��劙�jv�~�X�Bn���u���	!~�+��nv�,�	�/`�#����c����C䯷}��-��� a�l������:Qy��� T��<d�Y�I�p�ש��H��*���Ù�<[��%��8m@��;���~G���~ҡ���M�J��|1��Y����K�&�>����i7<�Fv�nj��SZ)N��2�u�P΅Y�@mځed���PQ��t3���
b$������&iP+Q��u�P��5����T�}�`�0�J������^I�u��ˮHo"����	�{��/��BBI˃+1(럼����FkB��z�}tQ���d	��x.�+�^�	?N��̌5�i!7���>T� v��A�u�l�(/�X��԰�!�}'
9+�K2Py0�3�"��Q{�i9���yR�+�j�j���4?������*���K���N�&�� �	�/���;�=�)����� �7;�� {�f1Ɲ$�6v��R破���:��'Ǜ:���C�k~��Q0�P��ܘi��i�T�����Dч���Y�Kbh�k!�r���ws�fZ�݅�قf����)�[a��!�O�x�dͭS �e��s�����tMh�"{���:G3>6��Ho�L�U%�q�D_�0���b��
N�T�g;�w��m�F>��f�)e�D[��E-���3���;��C���nS�Q��r�1eD�T�-�ŭ��|����_�2y�f�KN$!�EJ���'��a��Kf(p����@��
�H|4[ş�OW�AWe�8�c���ƨ�6�(z���cAA>|��}L+�^�c���;b�b�5չ���d�*��}�����<�ՇA>l��F��F�̡@���S��R��g�������!u��g0������E�5�Cch�9ʋ+����:.RqO�������0]�o��*KO�OAL.��R������F�9�����ہX���h��C���׀��rk?�$��	i�%���2�^�ux���(��܌[�ֹ�t7+�P��P�����Fz��HVQ8)�v�d�>v�Ӭ2/,�X\�S�A1�zN��R�U�_��{�=x0S�TY��ns>�,��?֦��P�E7����̑�e�N�u>���N�4SKg��..�hz�W�>>���gV��B�^Z`�5�ʅ��m�)`<d�ݲɖ����y���i
��;YA��~,{}%�ˍ8��bŰ).Gӕ#� �.�:O�}eZL5I���}t�m�X4"h��K��m���Q���j�1L|W�V��0�v,��TT�;ʨ�^У +I�0�T :*�m*4>��W���A�p���#�p��?��JYF�����H��� E�*��\�=��,��i��U<�|��KD�f�}BBd�wqZ��岸��vTP�ϐ/��u׮�ٖ���)93v�K9�6��G2c��/�I�&H�m������nŘ`�.)���F��"�A�f�E*�F#}B��F�i�[z.��k��@������#7bߘ�FӢ,�M��Q�?�^�Ls��U�ב�t�<�,X[?�H�E^=���8�IR����fT�V�2���,��Ύ5शCh�m�r>���׋���Z^kE�'�œ���	(���~�|������oSSi�0�ATY�?q+a���'i�~)z���G6",�+���^��Hw�2H}�
o���
���.�:�G�D/�~#!ĞG�)�� ��7���w���=ْݛ�=�.�[^�\.'�p�O-��9̏�#��ά}���ϐ9���V���gF5�g�Z��$����I~yRb�?�N�8�m��|�ms��_i��G�
�v4�-Ss���+�>��r��h>�U ���
���`ɂ�6r��)T��E;Vܚ{��?C�}�A�Œ1��I:֖���{8GI���I7c��`������*_
D����m����~<�w6]wĭ�&��:�ZH�h�0_
uy�-�6h���P�?�S�B\5ac��;��n���g� c�M�?b��7A�U�'�KܼS���VE4�|t�\�g�V5��1�@�=k�����ց@/���]���_�d���/B�B��0�,�����A��h�h1�ivHW���=L�3f&:>�>��o�U�|o3e@�[�t�Ȯ�Vl"F���\��S��9ŎJX�����՝�We��^U֧�M0�mO|\���*ޠI�ӻo�#E��B3���{���3kc��C����0���+t�+މPĦ���i�WU�'xTE�3�q�m#��G���R�a	�l�EE�8̴ZX�SlFa�֠��&�*��n1|��\�eVK��qx��Lt$�v�$r�̿s/��c� ��ܶ��T�R�EJ�N�~_�<��6Uf��O��=��_p�� uɖ
sP�����S>���Z��
�'`�ƃ%��(O�'h#���>��KT	�׮� S hv���S����V�:�����������FT�B�*���K�	j:���h	��a�9��A��n��5T���O��X���d^о���[���,#]l;�I]
=N��e
����Rl�p��D��o�wd<��?N���.��S(Vs)�|�JTkƇ8R�2�d�+K�+���Om0�|
��5K��6��$���W\���R�� ���=��%v��x7b�;�d�Qcd�I����|�6
PA�m"g����"!�W�E�of$�NU�\�5'--�㙵04���Wm��VTC�R�%�Ys@w��	ةu��Gd�. �nX�蠙Ь#v	kEؚ�36�9E���H�uK��k ��|��d�d_��\c�PH'�aU�����\�G����e�a4lS�$���Wd��'�?�G[X��>8czl1:���ۤ��R�����ܬ5N�>P5���o�0�w���m.�T���"&�JTW��j8]�A�|e�_���;Yt�t��4�l��хLc;���(���t=�kcZ�HI�M���絟΍[s��	M�B��d'kf�}�bXH��n�@>���K�&�m4OEx�+QҮ�Q}:6vUv?��?�mI�Oɀ�?���"�%�\���ȀA�Ui~e��� ���8P���T䈛�8�qΎP���G�5�� ?feIC�������YN�ƾ��3�A�`A�=n�� � �*�h�R5�_��K����g����{�1�`2�b�8����ؿ��"j��������F�:�����e1���9�/�i&3U�!,�Q�֌z�1Ԇ~�+ge3h<���J�4�#Cp��ZQ���ހY��{>05��% �>�h�y�o�fWn�[�قBcG�/:��c �s��*J�0k2�1����E�v�Ö���ا[���G��MhY������	e��E<�/����t�@�z=Ԋ�q��r�����ʎww���;vp*�$$[�b[�O�[7	�(Ģ*�'#�'����)�|�9|��zn;�,��"=RF��m��� ���W�8����lP�Ԍ��/u�oEtVՃ�;�].�%Z�@}D�?��pL ���^s���7����ܡ�[���hXt��Qt||)T�������r.[�UK�RQ��4RꯜL�o�""���{�:�ƪ����B/ck�CJ���)��3? (o��)�?���2�,��[���ƂY��Rk2��i UD��aG�_V)n.P4��f߉md-�}nj�5.�&к{��^� ��`l �e/k~��Niʡb�Z;�CO�*�GN�ʙ=�,��G��j��F�(�|x�^E")��d�b�Bɍޣ.<�A��ي^R恊�R`'3��<_J6xH��;�4y�l�>C ��_��RT�W
�L5����;��`�5��+��]P��r�#r����HH���^?��)��ƺ*}��8�	����i��� m����7j ��'��S�I��8����S>���x��e���-c����G�-.�t�i�P0���ɽ �b8��p-�/�NSҌ�X8hJTd;�u�P&���N
�Ł��7�Y��n¯�ʹ�����Ӽ�*0Uw>�� �IA�uX�O��j�(Ն;[s�x�硇��|�{���?crLc��j�iU��t�����0���ϥ����	m30}A3��
�St�+j4끹�a5I!�Ġы<E���Y��,vJ6O�Jo�lǰb+�w$� 7�@�����B��JB����*Ka$������fダ6������jx�{cf+����񓟤eA�T1`.�*�\�M�S�����c8I���)vw9���e�m�uX���o\L�М~(sR�l�Ǫ`~Jn
U���N��2.�Y�	��9�`��-�gxU~'  �kSl�%�q�l����L1���51�s1.�^�)O^�����L�0<�wV!��j��&�Y���V<� �"n9 *�=a�7M���Oc/���!(��b"_��m����� H�˞i�ő�Ŀ��F1�i@қ`����mw�3�?��,�b쥖lZ�Y��N1ݝ�G���#�?��tܩA1��U�BѶ�^J]�F�x_%㘲s&e�����^�kD+��`�Jr�ϒ�lC6a��)�w6�CF���G��*�h�Ip�%�Yp*�<�1l�D�i����{��v1��m ۰59?�i*��#�-=���ǹ�vA	�	�����+6�r��^�,�$28�at��Z�[F�E��5<�=t�v#�cL�/w/J���v�A���M�}J"j�s�Ur������ ��1P��8���f칋d�7�ch7�����e9
���ܲD���i�_c9.bm�@fc1�S���|��S����bT�D�$p�gc��6D�!�P�����|��/0	�w�#��O3$f�ʠ��o�*����I��c�^�8����u�VX#d a�	�������R��O�k�vzF�~�'��Y�PnV�\)�Լ���!��c3�g���}��J6���֮}]d�[�&=�<�c1�?�d����}�b�ȁƝ+C2���:��8�TW?����Ѷ��;��`��&/�����܄6~x9Z8kS�ޏ���4����i���+�˴��|N�Y�ܒjY�.����އ� ��#O�*�ZlH*��P熦L)�M.�� �w��t�9�f ���b!e�c���)-�V�-�F!	Z�y�S� -闚5O�q���>'-U�{���z)�5����'��q���â��U�-:ӟ�pޕ�x��SGNé֫������]���q��.o^+�@DR(=T��!DQcB�sD�D=hl�ɦo8�r?�:���I�hC�9�`�����Fg�\@n���n ^��MkH��6F�Z���
�k�xGT��%����?��ȼ�ŐD�Y�63Qf�=X�О�{KO"��l]^d�V۶�>��Φ� (��V�Ե]�ؙeD?�[G�A������s�	e�ΕD���S_��=�կ{$�Ъ�U!'������PL���������BjV�X��P�K��XL�������w��N�7�s_�9�jJ�����\8 �l�Lo� ��8�ck'#�0b����3w3���G�Sre����ҧ?��Z	�L�e8�����i�	����!��Œ�:���Ө��<erM+�շ�*���\���$�� %���WG�i��!s��-��������@�>���d�ބ%�҄���.�O�v3�t�޳�QCQ�T4!�v�R�
T�2�I�p�B3gO bkH�|2ב��@��q�C�D��.҂a,���}��P��@��8"�L��%`�^�����;|?�^�#�Eds���"K`��	G�9�6���8��n洶<�TP�#��Rl�%Kl|�;mp՞T|�pSVw�7���i8�S�3ݴy�8~au|�=�$~�!�8#��&M��O���TbP����_��T9�4�K�X�&�P��F�m�K% ��3�K5���X�~^e���K9v��,,��P�?:�bI�騨{��oK�����2����l��C��E+`�����J�/�)���M�$�G�5���V��]�\���jz�؝��z;߷�N�OG��8#�{l	�D��*U��$�����ګ������)8�Z~�xk�*)�Ë�W,yh��@$�j����2i���=BFV���eM�}t�=?%ژ�`�)������`I�"��x��G)m2]܋�^�!�EE��ԉ��b<�䍆S5v����:L�ɵ�~j��'���3-�T^��x�+wPig;������=�&��@��	x��Y5ï�l�t���(B�!\��"9�� "��M�/�_�K-�1��Cl�%ǋzTt�U}X�7j�ܩ��$oR���bM�n�z��I�V� �kUb֩陸�Ε����%
���j���f�������(��P�-�;k0�`�$$��6���F>���b>=���;%-s����:�ž�{D@�'gMΨwbة0�D�=.��K�Ga��ħ�lV�'����:��y�c0f(9�^���?�x���o���'��$�����'��z�2,�@� �^q"�� �0�h���84E��I��qj����(;����$`�y	�-�u���t��U�
D��|Δ�ӱc��ˑ� �`�UrS�N Y�8S�d����2����4s�B
�(�oh����0��Xc>	M���u0	q��p8��^�z,�]��U��:�%q��$�mZ�W��pkq^��� Q�/Q���	����J��:�X#&�t�y1Y�O�����1�)�w�v�BR�W9��D�)��.���|M��V�}^S)�S@폌�v,��i����R��nLh��,�4�D�98M6�έ����EM����V��H�>��it>qo�Q�������,wyx�Pb��|8!�k=�j��{���n�NI��ud�Z�Kk^E��ͳW4
��ͻB�s���l��Pv-c�%8���y��zh��X��!��7�Ou -Aw�o�ɯ$�����.+g�2O�!���87p�+n;l��~���í�˹��Ϛ{08���o6J�RHG�M7��y|�{��_�M��+�OF�E�O��r�geܩ	�Wݠ��t�3��hazY7�I4�{�h
�W�l�9�Adg����o���q�'��(�
d7�ū�{��F�a��?�7�RC�A�bڄ���f�@I����s��p��e��xg�>n�f	�HPP�&��z|���QX
��
i��QBD������>�EX���X���\������)�ە�~v}�Tɀ5"G����+w�Dm�&��e�K�{��>.���5�ms
H8^�0��\�]M �!黃t�iy\�#M����>ɍ-�\�#4�<Ű\a~����R�!w*km�A��^erеn�t����xl�������	��\����p�`Lv32��Z�'���)����������V�gq%��]U��,�(u�-̝��P۞x� j�u���Rb�?�b܀!�	��/�j`��aE�Y$F��t��Oak-�m��l^�]Sؤ2��f�E9h������n�0"3(�{S���&�s��Q������^�M�ԛ�K�_#g+�Z��v�B���I�5D!QHN�M{@�,��H�iZ�����8���[��h�[^Ml}!a�I���4��&R�����廽��0���b4��t�RȬ���Ef�۩�Y�����5z#����! �"YS�A���b�M6��r֎��c�-���Z�>�!Cؽ�-���Z^X��~n�~�����D��R����BK�!��Co�l��w���@�jr2�� ah⪱�z<7\�ׯ��I)�o���z���m{¤,��������v���*�����4���[����4�?����O���ႆ�����$@�ɓ�i�q�[I��*��~��_:���V쒼�K{4L釧�W�pb}�$�@�,�	���o���%"VE>rV�gT�/Z9�oh��1Ꮎ?78�Gݧ������}��^�l�̖0$e��;���`d�C�~�Up�I�צ���86���'A�s&�)�l��ma���#^��[�ЫD���Gr�`���s+a��T����>��x����5H>h#̽2�!��t�-�s֘���J'~9N�J�XCө�[h�f�ð�l���� ���v�.;��Ӯlp�?H�E�D�O#^�$��9�.M��N�����/�/��E���B=��t~��c��X�TT�H�����K�jGz��6<�VE`���g7���e:�Y�ߟ��~��'=��艺X�Mz��&��u(�$����9;����Gv���m��F��Kf�QK���� ��p���:�����e��Q�J�6H��ݻ� ����Y��6��22�	�����@��y���6��-�_��q�LU.O�=��yH�u���KFt���8�N��&�[$��pQ�~,�u����8��ŭ�LW�΅�J�i�9�z�˜.�z/^	�A+tjj&Nv�י��I��F �G�\Ȳ�.M;�=��}{� ��G�	�&@�%��o����8p�c~GQ&`��C����|�)�!��n&�5,�cE�g�	0FX!���<W,�ǿεߞ���� �';ge��3?��ϕ������ �{��,�&�1� .Lw�F"ʰ�L�R��j�b�0�bG`ƻ(���'`H� ?� �}KEl��.��ݙ��q38����jE��CYj�Ѽ�oJ:^�K���^��9����@��_Du��w���������-	b�fu��\�_��*-��{A`t��$a]i_R��pǊ#F����?�e��~�ɞ�{�<��j�}S��Z�"�-&���~���8;�!JdJ�S��g����q��#&�ef����8�dG�͢��4�EeɃ1�w {	�[�5��ƢaM�|�I]y����B��G=5a�\��L�5���)J�������|�U+�Oc�K�/� � R*�fU�;��T}MK������(]2�4�M-+Z��Q��M�g��p��*��ېy�h�_�lT�)Ф[紸ĩu�9� ��]FO��s�}[�&�Wa����#��pnW��ٿI��H� ����fL8a�x��?[���B�	f�
ʯ��P�L\�H# U*��o�o�Uine}TE���4m�	F�[r�����vީ ��� y[�����e��io�<T���7���P�-s�����MRَM h��]�N�s��G��̡<��XT�l>�)�a���^M��,�`�lI���1���<Ӂ9U}�^�2J"�M8��y<e��t�[��eX��e��������c�G�.��,G�1��ԍ�Y����'�%��F�Ö��.qd�V�8�Cvj��sI�y��l|����
���G��GHh���]�Fc�x�Ӌ�^	�]_�5�*9�rH��$�88!lC�<)�^��߰��8��b(��i!��=������\_ЄGR��l�áe(�}ڍ
R�`��I"��.En���}9�YZ[b?��۠oz��Z$Q1ES0��/��`<�3"�S���j��-�h6[7�����rB�l���-)�Q�cEs1�B���4�Ys��տzph����p��=�.s<�9��xx�
o����nL����d	)B|J�y���#IO�K����T\a�ę����Z�)��˟!�����&NQ8eMh�l�ƚ���(B��t&m�������6���C�D�{;)�%�K�HO)�n`;���F��f�kj���n�iN���E��b���i-����y��I-y��H�O�6V���;c&�D�8��q�OD���$����RJQ�6*cڌ��5;����ѣKr�ky�V&cy��]��c4͍�Qɂ\	�j��G?��u�2/�.Nz����XP�=��&^W�9�TcT�p�	�j�/G�<Ҩn� � �R�,�P���_͐���ȷһ�t��5k�e���DwR�3�<��TK~9�D�Kjn����P͞�^�S:Z����c�f�u)�0;F/7ܬ�٭}��ÛAR�����4��$�9�YL�ŖBy6}G�?�
I�sl"�2t�����?��z�0�W�L�_��c
��(��={[P�e����j��U+����v�~ih?H�(j��X1��� ��� |���Bآ��fV��Rՙ'h��B��3�Շ��ؠ�%����p!}���`��CG�Y�9�����!�z0'�$�-�(�]�&�X��)�S�և�x�]����	�G��,�;��W�.]�l�Eڪ�{K�+���G��=xό����!��.v.�3KaS�i�%�������:=w%de9*�+�9�B�3�N:���f?���&ͳK*N�-LW���>s*v،"`���q�$���E����Ol�q�4���Ϫ�6���5��T�0�?�3�����l�"X,i�>�a#_���9����k��=�Cc��"�Y�i�m}ѳ��QB ��_�0ѝ8۰C3�TW���_��&
C��匾���b{�|��qYP9��<�cmE������\��"�kF�|��F��m����Ƹ�;���I�nH�D��XeP�k��*J͸;�/�`E4 �s�N �@+�P��^���cy)��xK4�����
;���S��ł�LΨ��T9�xn�B�;���ڻ�z���KxFtU���I���J�E����ɵ���v�}g�Jăy�<7�1~:�6ͨu�����C�[�{
�.���P/�s�|�
�`eum�}{�B��<��{º>\X�*�Gn\�����$7��kc�|��<�E8��o{���ؙ���6P���د����p�{�H��ͺ���)�`��Iy�}~P��Z�(���"��tx��b�6!VR��Ԗ�\�.���G
�f�`�3�|�B�-����QP�r]��Y��~�	>m�h�i5��h�����,�la=�}��8c���׌JEf� 7g3�� Ul��H�K��9j4�UL�فh
;��r*�aU4����L�p�1��8!���H(F��,��|��6*n�ž�aw���Xí��4��)JZ `���߮��������)��+/��s��OӁgsNq�K	.�uS�m�H~�wDGd{ `�\�HW�G�̏�a@�(�FL�]B�h@���ԣB�;�]l��B��۳�0O��J)��K��/���{��N�3
�l�лX��oP�����:p	��Q-��LE!����&Ԝ�dR�0�~��ƿ;;�yL߹n��5l8��ʩ�`��e��b�h�a��{�;K�����B�����/V�ǛA�
\�;mN�:���4B��u�`N^�'���ĩ�򻷃��w��g����M��C�7��+r9�����.�O��%Yl��re+w��=���t�JoQy荼Ȓ���W�|�'*�S�~8m1h4(����n������ Ȥ�е��ڗ,5����:0�"y�c�"	��χDF<�sb��&Nܭ�r��6�r4,�tu���ߺ:#Z�>)9��b���j�K�}���}�;�W`�؉y�q�u��"�ϫm� ��ytG
�x�Hj4���~�g�K�wm�p�:���2a�,r��0i�!���o�BV�;%x?=�����;�|A�+,�+5�p�3pHf{���u�&�{2<;��g���0<K�%��c�f����F���#'kΕ�0v"����C��P}	~G�`R%,������[��i`a���a3�8^�O
�����pΐM��=��>��pE���ܱ�"W���>�Vz��^�{�N_�gW,T{m]�w��el�U7��q�w!����n�e�ܼv���b�
�^u}�S}��QeÚ�b�T��`���8�����H�ѭ��P��@�I �5��qV��@��+*�>|N�
!��.q�g>L��<���I��.�3�"���{���M3��ԉ��-���(-7Lʉv���v�/��L��߇L��bHP�@Dמ0譮�)��RJ)�"��f��C����xHd~����)K�����H7F?��m'��k�%�6�J7]0�����QF�ZP<�*��˽%w�l�'�]�#��M�`�������g�p��$�mP�[q@y��N7T���5�{*���	J8z
�D��(\)�M�|�힩��,���b�z�`���FݨLr�+�eF8C>'s5�_�ZR~Vu�QCTf�H��y�|��b��J���?=��f�|Ţ�JzP��u�MTD�A�܌=vr�h3��feo2�;-���Y���s����`w�7����|��1i��%���<�4�e�u=7�!�󸚔��,��*j!hM��_e$g��+�@��c2xčwW��%��{���"�x<|�wj�5�å��Y�-'kF��U,Ɔ#>Rp�;��8R���eLL]XK�?�� �Ta��wA�{�>Ȩ�#o��Z?dX���C�-����O#�kd�;9�6��vFwƤ\�oу����_�hD[*c��'�ř�Cq�{������:$��oԝ���̋�0��ȅ�?!?h��Dlԩx+ը<?�A�!(r�(�L��(&�X�1U�:O�"�Ӽ�d��H�2i�a��q�����v%Kz.��^��CHR,�+���p�gqĿ~�
���Y���֮���Ҫ��彔T)5ʩ��<r��Ӫ����ϰanpM�b����Jr�~U��ېW����E/�|_h�eU½�oD��D'�7��p����]-�}��LM5��0~'��㑜�E-�.���dp7�'y�,� f��@��ϾZR�]YO�j���� �>W�9�R��;ߤ��Vy�}&e������?f���1�D���4 ��t]����h�m���SYk�����>5��\�	F�0�*s�6_�â%V����V�袂a��UrQQ�^���$q9 �A�Q_d�y��A����n>��K�*֞}�x�+ U1i�<��-n):�V͈o$mè��~��ѿmP��6���sQ?�_q��u����I����4^�߁]��K-����_��s�`���`5���46`l%�F���/�>��l��z���ؓ8�WVHx~cݔ#ӉS@������d5��HZ�n V��){��f�`�&*�|G��n!;��*�<�B����k��YD�_�4-��hȱ�}�9pO=-���r���\Q���CVF�W�yb��G�	>έ��`�@&����hȊA�{tN0/��^�����#�L�@�Ki��N��,;.|)��v s���Ȇ��UU�kE+�]T�����W�n|����*+�S�c���&6g�c*=����x�-ܗ��\Q��~���w����K��V��u�Q�=s8���M�:�[&��B�ԚU��EЮP�õ�K���;�T��	0�|�L�x�x}��K}� sg��v��	(㊲k�M�)��O;�پ*�p@�r�$S��8%n3ت�6^@pT��~�R��}%tCipP�G��g�
|�U��:��0Q�|\@�/��m��I~�]���;�D��[u���5�f�(��}ɨ� p�H��LF�&����a��;t��V=������~�0������Ƙ dX��.yk` ݩ%�DY��a�T�8�}Ŏ�n*�Qf�8��LE�G��{�0��%7k�0�����t�WN�l�76*�������R���%��+��qUjF��{F��F��N�e����y����טA.3���d@X&�Ae���D)���BMkwugU��i\���>@��q|0��E�#d"	5�ӑ0���aԫ� �@���f��C"�'�p���KѮڢ6��!�_nۢ�0E�!��)}�PY�5��-멞P����3�V�1��u�}��Sِ��K������ֵ[E�Y~yP�� ��l�A�	��h5������@J�rD���=1�JG���^��k����N+�/�xU�$0��,��/�����r�vM�D�nG�C������>ܼLAo�`��]��&��-�\Zxe�6�:��ף<�@rK�4~65:�+���8rJ�~�Y��XY3���f�����\��_�{�^쬧.�^g�STs$<��)x]�4�5��J7���g�������z� �IJfk����X߄�31�1*G斓nߢ����x���X��`���$Y���0�$�O���-L��E�7[�5v��?�aK@�$����NM�j>�� _�R�
ݹi֤`�T�dd�7~mbo�U|�A���cG�q�^�Ӽ8���ҿ��?����g��9����RBP�
d���_�؝3���eߋNi�$$��O��S$��s�h��.��]������ ΔV�)���`$nE�S�����"+��G�����Z�_��(cN8�t�=�%�U\ -�n�wW;��/�pw��2���	���/JD92�~M��N����ƶ�AO�g�$N-ðk{���~s_�%af 6�aSɻc�~���<FR�U�ԋ�93ӣ�FSz)�v�Z{0c�^}shc�}5]x������f�\%8�bQ�A�mTgn�1�m'*gq��hR;�y�SC��Hqo�i@"rw�Ą�ZD�	���;��V��\�!�1��5]��tؖ*h�_����P&7jh'B�U*7�&���h�+��Mw)Rq�x���Q�� e(�~�(HD��ք����88����b��M��6-�b\�]+��O�����=���49eڱr<^*aw���j�'�3�]Yp�� OQ0��mᐬ��f��Mt�#��ԍ��4Bʺ�2�hռ�^�擆G���w�7�Zi9�Yc�q����/�K��t �i� |�پ�"�3��|y8���ǭ��m�O�&�Ѫ]��%O����j~gW?B#�H*v^}2�ʧ����^�[��~T�9��[������칰����M�if�-UΗѬo�K�.��oG�i�,$LR|�����V��g%T��a���l.S�_oxϧ�t?y���pj�J_-��0�O����tW
�E�a�!hk���N�t��*ǎfkD]��rG�� rl�L\-`��ξ��Jٜ:W�;Q�3YT�(���
��piI�AȌj��N��4X^���G�@3�?�!���Q-<C�V��N޳B�����4�"Ao�N������Q+�0�c
��b?�B���<��Z5��i�3T�Q:y�Ds���b�F��}CR��Ř߱�h�.�e��l����F�������h�+�M9�]�ds��������t�}��nz��a��n,�ҿ��g�8R�7n��a����V��@��'eSP ��|����_I��m�=B�
�]l��`X�Dؽ�X�(Gi��L+w�Z�����/w:�v����C��E�glq]�
)��f	����%�,�� �7L��"@C����2V_�`�`YRW6q�{;��D|�+��^"�Ͻ����f�V�$�@Wa�B H�׹CXFS�[ �]Ζ��&����uB6F-@�����	��Y�
j\�!�z��`T{�FN�hI��b�t�ni�+y�1+�������]wBH����x���X��`�ps����̔J���o�A%����F
KlϘvfU�)ڒxT	Ǟa�d���9�,)�2�L���d́��� I�A P(֔8+���[K����٠�>V�ĳZrP�V ρ�@�[�!�B�8���yZ���A��b�d0u��g��Qjr����ޯڛ�>��8W��n��F����!�h%8�s_�����ϠFB�[0d�w|0�I�#��oFxJ�#�k���G� �wS+�rEl��D �!Ѱ�����<� p����(��4K�ch3ְ��$@�QE�h���7l��+ t��O��n�];k�@o��-<~���;�������L���a��B��9H�sgr,$��m=��t7���OJ-�QZ�|x���O���f��k�`���(���]�2���w)�h�	ϸ��c�( ���x)\�[�ĕ6b/��4�j7o�7k�N<>[8(��>+Mi���*�)W+�aw���]��"56LǻGL���3��+Y�d��F��mu��U�[����r���=l�Fv�6�L��h��֞N�Ld̪[z7��R֭�ȼ9T4�@����n���'����6����W��v���p;�pf� ����4�^q��;Nǖt��wO8��.pbVm]yW���T��.:���k�x����O���Mhe�I~�6�Z�z�_�m�f���%6��8�a����H'zE#_^��H��Z�.�?^�i������,��T����g������T��ؠ�!j�'��Z���[��ss�B�PE���Qó�f���.��Bj�rxÃ��F����x�i97Ri�񾲯�.����}ۨ�_N_��{�_Q��f��<u�e����cRմ���{]��vű���4ܟ�(K�,�Ha����;�iثgo�Zтk�v�������6RRF���EB�\��O(�T������7ݴ�̏�` ��z�n�x��Y�v���	!.�_���g��?���hI1�A��kzD����w���;��ߴ7`�k�C��ǵ�L��XDP��p��ꔔ�P��¤a�i��j��c$���@"S<ɜzc�̭y����2���7�e�?����q�������k!����L��[m����~{�]x�6ƣ��-�}�j��Zp^)5�C�>��]ZJ0nf��Wdg��9�L��c����qĪ��wl�h�n��*/���P�z[-~z�&@1�f���{�M�㉱SiD�Rض%����{-Ի^�V"�'�ga7�Di=ö��Q�^���pnV�5X��|R��B�tq��imm�+14�X� @eZ �M�AD*g�j-���$��C���|�����ގ��w�ՋEk�w�v?qi6b�ɝ�!���z\L.*?"���h�
.��4�I����D[�E�Gs�ܦ� ���=7� �>v��M|c�@#����+S�t�#�����М�o�h�C�\������ߊQ
3~~y�ݥ�]�����)^������uB'0�[6aa�y�r��1�R��h�,��*l����6�q	�����Iٲ�g����5�P��/;��@˕kM�o �1��)���7Z� ���ѹNP��������y��y�����e6$C�I�V� ���f;�h{�b�:ƕr�:tIϒ�	�ɟ_~Ͼ6��7q��@��22Di7�t�X�����_��yV���V��l	d���"�o\vA�;Z4�4�~]��v�i���R"!F"~���������\>)y+�I;:!�U�;����Av�|�����}�7e˝�K�rؼ#x"���ZclL#aW �r����P�~K�Q�X�1C8A,�űI5�R�/���?�Bu��+������s?��~ �뎢��#;{j���&� b���<ނu%�1q�z���<���5~՝J<p{���ܺE��m='c[�HW�m�ɶ�	�؈�4����r���g�1/�[��%���������M�y
u����~T�#ņq-�����|�-LgA.j� <���Z�w�׾���<���S�������9�"�޼��UC���6��ph؍�����-��;�ф���:[N�3���G�j�e��EC�ԶS��S�7�������K��w0��_����y_�!!���f�N�۟��Ǥ����M?5{�A9����B~���0e4�c|v����)�Q򔮜��勞�����gZ��F,��|�Qow���90����@&���Kf�	V�컀ϔ���U�w�|ڏ�	���VM�A��K\�ye=e�ȇ}:9/�Q�<2�e@ÈS��ڶ���DH�	/�]��W�6;�*��=����"������3Yu�ɉl�n�ޔa9W7A�7*���1�3�\GN��V����i+p�bk�����7�ro���mOk� ��z���r�ȩ;{3%��Y�K�fiBx3UwIGFH%��]*:��E+Hap�$�;��.�ê��������_P��T4��B��ȇe�,���+�Yrۑ����P�Z�W�$s<ᥩ_�WD.I
+ŷ1��9��^��&Ud��Il����/�)� E��2�v4��3n|��P�8L�/�� i�vW`m��.P��#d^F��u�G��b."Ψ.�^ ����H<���T��	��m_A[~=Djk���f�d��c9�����O�ѣr|��n7ӂ��2y)X'F�:�=H�<w���n�
���^5M�G��\�-j���+������5@@0�keM�m"�X%���k���t9�=�6�LET�G=B���&?@	'��/��'��Ɗ�B�4��2��ݵ �T�hQ�v0| ˡ�%ҳ Aw�fv���@kd��ؐ5�:̒�y2e�0�	밤�>��$��#����1m�u�Km����q1"�e�	Di�g�]qM��u�\�F�a��ῴGKp���,+S��r�X<��}�S���)l
����+��R�r9��@�<���ۙ1:ၻPͬS�Δ8��Q6L��ef-��Z��~[#^�_�����/(�l�=��ۚΦ��7���i�
:X�3x9q�r�t.��q=��X����7�� ���܇;��v~�ʝ�C`��rQ���X�����$U��N7S5d��bT��J�xOCl�sJZ��{�wV�����p�,�����-s����Tk�ɺ������Vޙo�R�Ε(1�4�a��f�`�����p���й��{q�O��b�𼠯L�5@>�%�N�hQ!�M,)fTjb�O!$����0��6w��"�d�<�,{#���QufL��S,w���c���Xl�<7Oڦ+�_ �����&��l�QG{]`�z�iFKk�x������F �ۖ�)^��+��ᒁ:�ж�H�wx����tŚ?O��8U��T7נ&Blb{ś尩S.�v��h8�%4Y�����;A�I ��������4����P���A���͌P9�;[0���W,Z/�%F"��B�����=W��C��T�0�I&��fZ	����M1w)�Hߣ,hL�K�3Ķ�K?%���]u�u�i	n�����hѳ�m���:�l3�J�3�_K~$a+s��\C�'���!?�C'2Q�B�W��IV-喝���r"���6�o�4}ʨ�%���K�M~|���!�p1�~4��\{q�<�(Ig4eL,nO���b���d{D�~�ڱ�m�3=&�H5�I;j����rk#��[�h�A�����[	)P1u�&�V�>�¿��)�������;���v�9���8�����P�u����'�J�{C\/��Zز��.Wz�����ݗ�[�O,1�r�ƱΧ�2JF@���LKk\:�t�寺���;I���4�!����Yʢn�8`W�*�P��!�L.�����Q�3HL	��]����R��Ӱ��v�XC3�<�Z �,��u�߯�3��/Q�JEG���%&��`:�� ��׏R{Z�<Մ�j��q��g#@��:Q��h�$u��ELF�`��"J�G&���2c40�A�a����h����o�w���"���%�_p��2�g]X�[�����1�؂C��<�y�o@z�p�%�J�G9���r�B��'*#A��f4���KQ�l�[<��{�qg+�ϊ���Xo�Y����]��;�O�|������t��~�C!�	����.�>�꼉k�^>�Wh����}�	=-��K� ��+����qr�)��ѵ����^(��[�������h�l�4@�^{0?���y�ޚ_�����֔{
l�돘�HG���K��6�����i�
&�p�tWB�j�P�ׯn��z���
��qu���Ԏ�+���Y��~����[�ѭ�wC�N��v�ʊ�0r���"y���m_���ɘ!��1X;�o��7���6X*dN$����^�
���ԛЃ��k�ȿ!��hް�v�8۽�dV�<;��������{.�M8�@���V&:�
���H͹���0d�����X*C����/�K�h�Ɏ��s�;!�U��%ѽ%H�)�v�,"ذx��;��{�
�4
�o"Y�OwV��\|�
���Lq\w�����5KA4�
�qVu��*@�JTt3~�Y�7�ۍFϭ7�Uy�j���`�ble��Zy�1 ���H�X�=y+����*>Z78�R��.�D�MT�i�G��-iQ���sH�T�țV;Z%
�+�V�H�՝�V�I*3y!Nl�MT���:�r���*�oR�%+O_���/k����YǏ��R��X���d+�-��a����2�B�J�H�]��yh�L��ɟ�FZD�'���|/XҒga�gJ�ćs	���P�S!�=�R��̿n�uQ�\������g}Un�az;Lxl� ��v��yS� �d2i	tttK9�����oo3ܾ�*.V�W@�6]�h���0���x�����C�����[�w�R�Ep�l��H������$�pH
#ӊ*ny���K��]��Z�Ta�z%0{8S�b�J�Yk6K�B:�[�a�a��>�	,�6�갩������Ƀ�`�����_U	�.�#r�h[NŌ�&�K
�V���L��0��,�{������Z�V����1o]��m
L��φ+uT���[z���۬���-�gX�ͅ����Ò�����Xʀ����}U6s���H�����-�+��$*wp�S�-g���Z'���"ag!����GJjpB'�K��DA(���
�����E���u3]�M=r��AAז���jK
`[�M�8��ն�L��xR�{(�3�i��6��}Iz>2̍-Եr�F�^����9���>�ms�[��ձ����HhKh]toj�=D�r�����H�:>��0+n���qMWNt�o��z��`��W�>ﭧ	����?1�k�VQ�_����D�ۥ��ғ�;��1�c2"Ճ��=;���?�m�R��V�!I�Ĩ��L�����7�A*ն�<i�c.�-ۣv|*�hD5"����V.40^�4��oyXE�$=�_	��v=���>�4yz�yT=���U���Щ�&�U���iB_��Y6/��V��3��&�b���h4��V�_�cW>���@ڊ ���)�"�%[86!61�g��\���+�R�z���/Q1)��l��;���,���}��?4��j�׺��@�ӸZ�s�8��9O=���&����-�$�J�����[��)4��x=+�$��r��4Kyh���������ï�$���������cT����m���C8�����3S��F��
Hr�:���S�YV�s�Rg�O����n��������p{[qT�|�-oTJai��p�/k�Ѡ(�{����{"s}#�����V ���DI��(o1:������5�RŞ �{�P�];�n�[ݔh�U�O2���g��{�v� ��Ա�Ql̸��\XN6�����^B�B���9�g<ñ��c�T|�kLӜ�1#A����$V�����I���r߬���5�[�K��5L����.\�-����C����Z���2Px�a�$vڣuъE�2����Ց��EX0EBrZs�bMf8ŭ6b
E��� 	[E�Òm�8}
��S�?���>d!���:�:dIH㘜f2~����^���pq�n@��3�V��8�}���%�?ɬJc[�u��������u?��xd!e��jW��Z�}N/3��Zχ=g�泍���~���\/Er�)e�䡘^�z���V�o���c�����5NpNB��]_?�o���`k��͍4�1��>E\�OL����T�B.��}�~t @n�}�"~u�ſ/[ɾl�r���i�"�E����o��������F&�NU������2n+�`(1]��,�i��|�?o��w�C��Cwo��a���3�2��ݗ���|U�C�m�i�P^>���Q����'��ɦ�=�M���m���a|y�"���?#�+�F�Y����{D�"�k�
�v�c�t�T�<�Fi;�2F�b
��_H�
(���ߨ�ٞ�k�7i~��~�����h�:9��D�&b_f�&�xM�~G������4g��6]����[k#�����{��P��m��7���œ����9뒌�RIv.��D!�ׇ��)%���I�����{J���B�\�ߔ��)R��,=���C&�h ~F�-{]�F�/]�g�󑻤T�ӿ}����eFQ��������{��Ĺ�{d�e��A+���_�6����^�A�UGE�ZU��Ph%1��B���`��>j7r��6>�{l�L�.���AF�.Q͉�}��b9ɡ�m R��Q/�%�X�8
��~,#�[�0�m���<1
"^镤�^h�����!���<�zF�����{��5���tNm�#B�8l����ߘ��U+���5�ck�{�-�`���$� ���� ��(X��"JS<��ӆE����3���u<OJ�oY����X���T�����_�i�Nv�J�o��0כ�[�{��M��7�\|z^Jɉ@Xua�5��୊�p7xGÊ��>ܚ��� ��2���|��AK�(��Y�l�xw���O�����Xj�s>�*�F˸��f��%���^K����G���(�6��!�vV%�P�kC�֡) LbM�d�Z�\��a�4B��EA֗@��r�_����uT��aI~f�r�O�t6��@z�W~��,���g���$�ye��L\��!g'����h$�Z�W�����ӌ�oޛ��|�wxNV�3�Ϗ	��{�����,��A��j��񐴟�J��Y���D*�ƶV������@ss�C��#/������rmHM������`+���P1Y���j���oƭ��Zs{���ΜF���7��13c,j�3� ���XmbG�y���f��Ϗc&,�	pX_���������Xy�N��i33
�Nٿp�\s��Ĥ�(�f���V$�V��p�<:"���6�	�ͤ`T���o'�i1EқVa�pi�+�t��^�Η���c"�c*�A�,s��H�^ެ�s����I *�+�����'�)!gLk�}[����K��Fzͮŷ�>��u�
��^H���r�6��Q�
�\38��,��)*h�2��*z{%��n�\�h�r�]�'p�����h�	�ۅʫ�G��@�	���&^�I:�kH�9,M�Mh�t�$��a��Mnx�Qe���nPf��6Q�0�_}P��z�7@ep3D�)�3�a�fL��e�?xt�P�3�x^�<V ��Va��(�O�D����*��b��SD��Y��R'[�;1�χRҡr~ �����Lm:������=U�E�����c'@(|ED�Dg3��z+���0{1�ŶՐ\�e�usm�4{���W��Xk|���sV9_~����Z<:.�q�"�K�U�Gv���K�jm�YS�zT������nR�ˎ߭PQv}J�@-Ă�m�΢�Q�>CM�yM��;[ As?6!>����~QI���0)j��Ӵ[X�<3�� �S����#N$f�����"<1��s�I1�8n�V/7��[&�ߒ� �h>B�GaiI��2Vٱ���v�	�qO������?������<n%���h���Wi��3'���2m�^�2p��O�<5���	��.�+�q��O3�Ȅ�a�aߴ��*D�x`�H^>�n /�� 5GW��2D!�,jY�� ��"�Q;rH�v�&�3.�4��l��
|W�G�2s\�5٣lɶ�a~�'���瘵B��,<7|&�E��?���lIYW˅Q}z֍R��B��f?o�k��`���[3\���W�W�Ѕ��}ރZ���X\�O ��sy*3d����3LQ_
�٘�?��ϰ��)��'��B�t�xi8��Ark�!���Vw*^��2�OJxGG��4��'�nH.����[�yꃟ:X8 �P|U/t����xsɋ���y�ٕd=5TUA/l8k[����e�h=��c�]݄jh$��:�S�<��Wa�)�7��2]8�_�!$A���j(�����4�8�S��@��pD��@�F��.L��&����jH��3���cW����9o�h�?I��
�)#��  ���Y�)X_XF��& L=��f�
n[�.F�Y=
�p����Z �,%�I�V���j��'�ֵ�*F,�Q���x�WTh�_;��C� Sr�fI��2N{r�F�Y��C����i1�C��ٙ�`�-�_��'$���Pl+�I�i�?�K���%n�[y� e4m|�	��o��Y�
*t_�pU�HV�Mgc-8��CЖ�g5�����/������Խ]�fP�����~���'��2�/ �	�P/M	��ǒ'%_�	��P��v�,�:q����nN"�k2��;��y�ã:��O������Z�,��A�Y�� ߖFs�C� pp���֜T�~q�d�Y0/��X�V.o� �)ty~Y䗿�a������N�z䬴	dV���}��$��U�_ՍO�t	�n��K��G��t)���T|]���׆J��U�#X̧�{�(���CRbݶ"_�Qɹ��F0���a���}��v����� ��
z2S9��C��	�E��v_O���TX�G�uzÇ�	K��Ŀ]+�n:	�N��w��)�{�x��l[Dp^�\����<��/#|W �<�����9~,�㺷��vv�"yI�޻/̖<eaR@ �|&=��п�-�|5��N);��*�͕�t�?wg㎸u����3�W�B��W�򈎹�!*���Oʑ���"��pb�wB�ym��� ���$�q<���{��{(������2����}��o�ʱ>���ӮJ���H�l��L�<�U"�iL����-�}X�J�r����9����ԗ�o>�1���A��S��|@�D
����ȓ��A�m��R !�h���f������i��Ϭ��7�c~ �`���i5J�xtQ�Ko�"@4�%Md�!����t�ZY��be������~b�m������kE�Π��}UA9>��	�p|�a��D{3�=
�C��s��"��:u];�#�U텉���Af2fM�#KY���c��U��o�ԻQ���8��Ax�O8�vĝ,��I�Nx\5��E��YE�.��#���4Ը�����ePZU�7�}�1h6�,ѼV���\Dh�?���~\�x�zkl��Y=(xgާ��������*�����ޘ� ~����/�h^�
p���a�m#Xȁ���~��a4��D�pXf�E$�m�$����A�y�����nFK���/p2Z .s[�4�M����	!	�S�C�U�`|2<sL6��!�oԐ�\�&�&��e��&��a
����u�
���#kRDQ�wJ2�����a���9�6��P�f$���s ,/����"�`�\�
TI�<sPʋ�`S"�hD�^7�{1���&��AUѹ~�4��Fڪ���@R�w�K����I�rll����l:��o_��П(n	�6Z�Qf����}u�J��mA����4e�W���w�A����	�8���C��/���3|�-6���"�Y��ysq{�V�l~n�L�ʇh#j��Ŭ������_��4�/&��"�	����T<�c�z\�}��h
I�!c�p��
Y�4>�Ul ,ZA%��{��n��e���°H���VT8�UR���ʜ�j����V�\6N��`z�T�.k3{7σ~_ȧN�S�s]ϙz�h�	��3,7��c��ú�Ng�b��
zsh�O/�:�]���I��7{����V��#5�P���yg!BcE�1��K7�S��cJQ��Uw�z�yl����;����� �\�+�-R��*�$�\���s���!�%yu��l�����W�� z>/�߭��� �����}��x>(���°�n�K�Y�n�ts-��ǵ��\�sުD7>�����>�f�������ߔ�ň�������4��є}}�����dNnm��\~����f�]������.&�Z	n����������r�ݾ�����w��9��ʺ�I�*Ls@?���_/I�J�	䫷����_��ր:�o�QUe��-e�~ZP&�Ҧ����|�{R����y˯HN��;x��Wh���RW�F( �3��^��}���Nཁ���R���+E��ljlP'eaT)��r"5,�LS|# (r�t�V�V1J�U�r�m�7�c����p�o�y�ګ�̂���(�� P[�H�G]�a:G簵­��ϲ���;��3���r*�A��L�mce��X|S��:A6+���4AL}lõ�]�d���F�4�Y�l�����G�n �F�>V��S��}�
_����m����LV�ǅ��?�.�[%�k��a�đji��ZU��M�ex)u�Km�f}3r���s�N����(��n�;�oG�z�'�`�c�u�颥ϜF!_�@�ƫ@�0��<;�?�������i�\�C	�[�FcK�M=���G-�]K3M��L�{5?�k���:b�g>� ��$D�,�W��Vh�[x���.��f��EM�+r'�GB��l<@�)��C�I�g�Z���� ��?�>�ϕ���:�E,d���R�<\�h�v>t���i�/��Z+��*JS�cG�l���9��-=7����,�~��N�̆��Z%��p�h8ߒ�<�: '�2ۤdP��71�<hcyl6�⎠Ѝ�^�	�k��F�^q�,��>=|�����6����8/-*ܹj��ք�0�����T䯸"G&���<�����G��,2(t��,��U�H�X��~҇�u"~4T�\B�m06�ph���ۦ�,N�s�˳��=��tI�D<�������c����'�Cv����1�������-k�,���};��&�kX$�ۏv�?o'�2���"?E8W���k�5�vOC�Oa�]}`*��e�gu�ydZ�4�����Au��6�G�K=Wo���}I	'��s=4ɷ�6*�5[���]IjC_ob�Fmp-��|��ib�i�n��6�?�H�k��,.(H�1qq�"@�g�G�c�"��\�y�P�o���J7��{�
�#�K`����`8:����}��� &f&���U�C�>	�t�`	���������,��(��1(��^�(�fŰ�GY��&���u]h,]���ۥ�+�����S��?e(����㽥�}��d��i���v�����ҹZ��v{��WY�*z6������'�|@އ��-��Lǣ*�v�lBa���S��7��ڷy��I��e�k�,3D��EG�gYAb��M	�A�#'�;�J�ݳt?8P_��Co�&���w��C�wtz1�(j�i$bB�Rf C�9���zJ�%��}�q�P˞;�M!�gz����w��&����h����c%�i��O-�NQ��癌�?�Z�!�a*�Ĩ�He ec�h6�	���bgΐ���}���#&	���:�'o�Κ��@i����iXד�x5̊0��%��r����� �8�����7��+�v�&�F?��N��i�D�����RfZ>g;����^���nZ с��]�,%�Ihݪ�s�G��xJЯ�A��4�n�����|�������
�k3���-�s������h�~mh����g���˫���j>����2�ߋ����ߢH��s���j��Mx� �w��Яϸ�����0:�@.uA([�����V�D��|����Ps�%h�ft�H�3�/GHt9&�V�$���E2��B ����Y���7"ƚ�zp�N�>n����߭ ���u�]m�,��a$��N�ϸX� �|��.�'�(��<���K����Xj'�Q<�Rhw����$}i:�s���+ ٰZl)��i,��p�/�.X��X���[�'ȫ�=�}�B LIz�+�p����W�b�qec0�-�*(q�}���z��0�HI��E��Bd-׵�=@�kM3�q� ��uL�c:7\f^�����igK-��_���wa�i�v�AJ�����%	f�X���H�`ƬUB�P|�g�����Ǻ�Db@4e���aر�yn�3�%h��٪�Z�J�on�i�7�f�
��њ֫�p�vF7=.��Hf9ܤG�A-�8r�/���4y���F��CDۅǫ_��F~���AȊ��n�����i
�N._�wL���O�b���E�^:��ߛ?(U�{;�~G���P<�����L��Yu�rN��J�:�xy%a3<͂)�O�.ܿ蹷c��m�g�S�4A_�;���@f�*[,�j� �x,D	��|�.*��p�����CBP��y��=wdjm��X�r-�S���{��L3�������m�'B!�ViN�25`'yRg�n�$g�a�����9`��u��ͅ1�YO ��uL�	���9�B,���H��"љ�f��Y�h�/)��1��b��G�-z��Q�����,A�Iɧ@�Z `��3��y)����� ��7W�.������0���T;�m/��Xq����2㺴=�@۰�ږ�Q�rW�q�m�ioׯ?#��
{x���e�t�F`u�����Z�3��Sg^������Ch�FYD{x$�T�¥U9�W��g�&�e�'��/:J���˼�A}�޶?�C[���W�^D��G�&�b��X���6����{�# s�\A�
	qh��{c�{B!0�N}���# {��@��賠깉Թ,�V=")�+�߃��u��-����sW�5(��3<w�d^2��l�1��;e�hdj5Ō����@'0WLp�S�J�FD��Y�M�YD{ �&J@Wn�W^��&���6�����&��.���YGvC*�=����2)Pρg$>F��ӬՒ	d�4�A)��j y".g��L�5f�u�����*�K�j`m�S�1��n��jB��굡C��$o@�D-���� d`�0|�6U���,������g��L�Ωt⟨.���d��1y���-sSfv����J�~ˊ"i˖�9��R���z�HkM`h�p�.�k��ɫ����Q�X���,���V�
Z�%7���Z�t�\ŭɐ_���$ ��t{Z�FRqe�Z��ߤ ��`%�sF9�cT�(*��-��B��Vx��U/�SC�o=��T6�sB]Q�~� CGx+����1�f��Vzc���@��4u�����7i��вUf-���ևH��R�zr
��7ώ�'�#����/G{S?�i�+�f4`��(�KF(@Vn��|����Ѵ�Z����}^��v~;|��<�KcJ�+��P)�N��C?V&a�k����H�[�ϓC�>W��Kj6��$��k��(����6#��:J1�_�6v�)u#à}N/8-������G�:r�KVe����I ,��t�[7Z�I�;��)G?M����?�5gi��I/?t��c�D/�WSr��ӑS l��<B�F$DY�O&�t����v	gZ^�"b]�}�lQ�U�C�A���:��;��h|��|6�uY�0�w�^n>�*(B��NV�*��WH-&�ll���a�+F7�+�����|�I���ck��|S�����<>ˬN��3�����l'��ﰘ��7��|9=���O@..��,�Z ���"��Ho�b�7%Bj����E#L��M����:�P�?����X�F�&��34��*
?���>����d@QF�8?���L�fU�E��y�q�Y��x�;1ݔ��w�BՕ����7��{�w^l<�5*"�o�ş��e�s�GB&�8Q���&1�vCPv2RN�tv�2�'���&&��ωt��{��Gs��Rbp�J���[�>�öT�N0ː���U��/c<���o�(��/�����d���=������A�0�ݹAԏ�=m��1��{j2NrmY#�sG�~Q~
��e2��m�4�����|6�` T�����3��4Ȫ��e��B�e�� Lb}r�9O ��Җ`�Z�7Q�ZX�Dl�޲����!ۄ�8�=3~���}W/�/�g\��)�J>����!wz����`D<Wsb&����Eջ����r�n��h�R`TN�@��{ʁo������,��n±;�-\�k�^��ճ�,ʾ0���+��Ql�^XeX��x7��ztub�Y~�9�v6����V��&���!�6F J��C�dVBBi�6��i��ewGhI�+u�Av[RoN��&h�e�.�ƺ(�;&&�L��e��u_x�
q�1�	�QL��$;Ư����h��~F�O�'Bmj��g����Pe)2QH#.]���K�N�E���Sz4	�OP��Ph���o���0Wҁ'@�sph���߭��r��t���i5��m��	�����2;��I�y� �6�f��Z�s1�.{(>s�\�CB�OY�G�_w��x��\Cfde��Gô��t b0�c�YV��5jG������9Ēx�iz��E�F�"![�J86|F�9�dx��thB�=�����x�P���-W$�z�� �[O��*I�[���t�@�6֜���o��j��Q�}+r�r�Y��;1�S���rlk��iȫ56�))�Eyā��G!�����d�M�.�Mh=V�Eaе^u���Z(�eC�=�����Fp7�^�ӼS�ʧ�f�^��ik�d
`.@�D���b�a�[��q~q�=Z�8'[Z�ϳ-�{3���/X�W�~[��*�1uI���-a�iϾ�@����p�ە
��{�����@9E���OwΊ�(X��=�z;�6��Aiq��1}l+��ȅP�]r�t��Ar��B�{�}�oސc�C��Y��c��a��<�Yi &����0U� �.ֹ�Wvs�dW�r���m0mˣ�� 	N^̨�)d���X��*k�x���VV��V���+�V珋<�wdy-�Fy`Y|�g�u���T��(��vda�/4{\���	x(2Yd��
{��ւ��k{�Ew��Q��1�y|8���v/M;*g]�+�����m���X�M���DN�^�x�	p�������Z��v/Q��®�8N����?/R����~��������aݡ�Pz��cdN��G�@xi�G*,��nzO�H:p�4��!�g�D�ydw�aRg?�W�)줤��`J>����W 6&oQװw�q���>[���(���ly{�[i���T+�TC��J����S�Y�Y���r8�J ����$9$jkV����_���l�^A��&ժ;���?�^?��5�NtkYީ�93�w��zսu�nn�������y��'3� kM���X�\AHz�y�����L��j+#
6�����?�N��U���쪸�xgl�r�0�$'³�����z<��1u&��9��Ĺ�����y칎HG����p6�Ч.ך?�Vᨶ����U�DR��\���y�ѣr7�ʍ�'h�ږl��ܞ�3;�\���m�0e�I��(d����4y��VȀ�R�w�=�G��ަVP�\����\�c�Ԛ��mih�Ν��57�9�'��s������l�&��6�_��R�I���r������0�1m��$t"5��AX�L��%TP�J�ś�3�U4��ʺF�]��c<�Q������:�����/]��'0K:���$t0:ʆ�#�������n]gScwy�
�xwj����i�J��,o�$Z�����z��X�狚Θŝ�
hRFA����ȼQx�ޅ(�o��ކn,a!2,ڑR��Zk*46Ă1��l��ᣚ�Q�!"T�.����~ϙ�a�ޢ�J���{�r���Ys��J��gT�Qy���]?�Ϗf���WH/�b-��D��E94s����:V�����}xر���.m�`���%RH<I��f 
�ߝ ����m��&;��#��x�k_�jN������1	6�B�f�q�n���+���э�����7���W��pi��4�� ��
��rH#"X�[�a�{�2��ڗ�'J�ͩwJPŮ��KT'�0�pfs4&hcD��@_�'�Y/��ob�*x|_:�@wlyD�{����vx������Zt|����Xn;�JC�/�e�d�T�;��j��y��oCU�y�Bg���>��UM�:d�>-w����G�rY��w�?��l��x��Ƈ�Q ܖqoN�ceF.c�m.JgmnD� �2�!q���V)���A�����lpS7FL��%^�X7����&8O���Ǎ������4Pݬ�� �;Ny-�\����������u+?��L�DzV�Tc'���B��
�;^����Fl�G�<Ѭ�ۍ��߀�X	P��8�������W�@۵���5����xjWm-&��y?- �������о�z�l�gLيn*��VRc��uR�Y4s-5�Ͽx %Fv=l~�l�w�JJ�A`*l��|�˺�<^�����i�LZ�+ڣT�Ĺ��
HT��ـ��:��(So��soѐ��_W��V*���m}�����z c���I�$�qy��\�����l�o��d/\ ����74BS�@sh�~0�.q&��a%�+�����Q����4XW�-1w�$z�ޟ!lU��tS�8���9��IT�V²�����Qe��jf�ڠf��3��D��h�����h�L,���-D��v��E��Wv\2]�(G�Ǎ�H���"�*"gx����	.}�L0�H� �΋����1M��EM�IK��;P�6�?��o�& <"�gAy4��
ɑhw��+�(��d� ���3G���ATI6Pf�doݽ�o��)먾��M@r��6��,6z�^9l1«�@�t%��<���t�y��	�|r�M��e����Z(g�������<1"[�$I9Ύ�����,H�x�"a�a;[`DyMō��6�p�+%Y�խ`����eѵA>�*�Cț���;�	3�q<̏`��Vi�~�k=Ǩ5�����N�<#a�j'W�3ҷBU�oW�����	�,���/^!�1�z��5#-�b<��Ȣ����?�&FY=AG�������ǧ^a�Ī��G��>��\��Ю����_�jۍ^]8=Q�����I��5��D�����Xh[�0��6$�E�S��_�cFDϦ��H�2A�}�k=��+o�ax�FA���oJ�+Hv�@�x�ބL�[�E�j��yX4̑q_�bkҌ'8����>n�F�ۜ*��3�v���@��\V�G@%Ι�W�d�;�bF��ߞ�E&�j'�h�miC�Q�~�v��pK�~�ܜ�@m~Dz��rN��>�K�QRl���5�R�1D�EnK}��F�^v���Y$����T݇˷��b*M; �3O��`ħ<؈#��7eLk�'s�"�;'�v;�L��45�k㜐R���f�@нLфZ����ɘ턄�������&����e��{�b�� ����̧�6�PN~��C1P �0g^4��#$����B�b���am{�T5S�&�N��	>>�RVn��#�ᖙ��\����w/�ʌg�����
�� y�C��[3��'�Ak�J���RZ
���Άz�Xox��ɲ���C�C�^V�/	?h�z�(��������I�Rs2��\Y۱���� Oĺ �pЫ�,-�U�_@��c�;'�SfD�[(��˅�����1L"����e�YCg2��&���|a�����}��j[x��c�R ��~t�*0����&�����B�e�hpI��P�e#�ޚ��hƞ�g�s�#��ﻐ��"�^�t=�6����6�3ty�T|`�+%ܧ'M���'Y�>߰�|����c����2�;�L��X"�4�=�V�أʺ6���)����7������sɪ�v���h���Ĕ���E������U��l{�
����4��2�BDQ�Nҫ����}s[�\�bx=�µ�v��Tí�$`����Ӡ�ρV�Id�ĝ��6r&&����5�,D�&����3���@����+L]B}�H� ��4�����:N#��X�{��ɱc�T���}����D(�^'�wdB����!U7|U[��5JI��f
�r�'�M���u�&�Mn��p�gC��z��~����w���ބ`�O��/1���ӡm��7�!Y*�$�z`��r�
5��r�a�u����~�y�u>�\�G���t9�� ���/(�;�fcp�5'��֢��1�G�G��������3��hDu(�d�k�K�.5��c�9�m��s���6����܍\���R�D����6o�R�Q�^[��{�X{9�ԭ���Q/S(J�n�Hkr��)0>��]�R��ܐlAW��hN� ?W7±u�t�m�)H�c!�P�Y��"�ὓ�D�]���Y�n,�|Ap(P�<H��9�QEo��Yyb9w%��5�3 �.	v՞�T���dd������Hg_��s������2M�u��8��1e~�eV,KzW7�%c����e�Ȁ�������C@8U���ah�&��僖��6�Z>��q�|q8R��<y��C`MI�*�]� ���'Ȑ4����@�g�O;zr��Y��B�Jj�>�F���Y#Ff�f�Uk����'�0�d��}u<�s��.ț��٬��G{�N�c�j�p�^xZK޾����-9��)�����kt�/�1�
�y~軒SN��뽁���/�C���ESF�	�<�}���  �*�|ݫD0
�7ʵ�)RA^Ejz��5 ���n^�Y*�椴Q�v�U��M��&t�:N$��7}��7I`T�&��2���+$bԦD��Z`w�z��i)(J�G�=j��Ǚ�4d�lyI�Q'og�X._���Z�"�>/E<��F~ڳ&��e�竛.��¶�b!��U��(!"����J�W>��Xڵ6=±hk'�B��f�h���\ ��g��R�iL�@�=�������-G˃3Y&	yw�'�F>q�Q�%��Z`{n���PxU�����_���&�L?g$�=u��%�S�[>�s�Z<+��ǒi	�����m�yG�=J��5����![�	���I!j.�t�В�����Db���d,����C����-�U�[���K�j�{2��B�@Eqs.��ao��K���!XV����p2k�s�]��+���(.����3lu����V�R��Ts�I=�U=skY����#3�U�<Y��^nI9A|_�]��{f�Y`(���ߑʽؐ�  �A>����w��	4��;��+�}�����9H�R�$����fI�&���z����7:������>&�����s�X�K��~�D)�s�`���=M_7Y�	����ݎ�C8]��OS]6��s�ܽL��eO��N��TI�G}I���M��fOǜ�֠(���Vߪ��nT�y�bn���j�R��x�Y�4�FԚ��m��+
d�'�{�~W=O6��5�m�(�COw��L�� ԊE>/3��r]��SA��x�!A�����T�-���FQ(�;��eO.Z[����S���ѕʵ~�<w�K�x�_���a�h�.�ֱZ$n��G��&Z�������Q�eF�,g�=z�w�f�/@V�K��A6��>�W?��� �O�n;�u�i�w<�ri95�	�P2�R�[�7�6�h�c��9m��)�a�>�E�ى'z�e�T�ȓ-@���)c�Q��i�5�u�?���+b1MK����1?�qdu��,�zvK��L���j�2�$����4��o�jH�-ٹ»�/~�ʶ7��o��)X�zj�E����\P��E�G��H��,�C#ւ�$>@�i)�+��e����>f�I�UO��Œ���E�x���mf�����ԯD�ɠ�lSz��p�jdFy���;i��t�} ���9IGO����~?�_U�ǋ%�3�r��ۀ~��@DS_���+�X"�@x^O���~ՕJ�o�_X�'�lN^54P\��'����Tεm!-�Rm���h+B$ςʐC�����z_��*Y0)�y��ت��A��[Uϑ���W���P���T��];ʰ�bd 3��}�+����N��I�����Åd��S\�/Jղ�e�/�ό�� Y���Q������3�	��@.�)�Q���=<�^n�����i��,ё߱j�+��>���j>��{����.�HWn�%R17��F���:P�,��ZKѹ(! �����S�2�Lz��{w���������w����^e�`?7_e��U��qWB��3K�� ���N�8gV�ڦ CJ/«��=6��rbQ���+ǔ�B*�L�����ہ��PՈS�4���8�[�߮�I+H|/=�d#�J��iѕ��K�����({���!��M��$���Ϣ��)��z�}�!8�e���)�{^|�+�Z�Ψ�*�����X���Յ$�u`ed�����G.{+E���#��PH�L�/�1`y�܊�DW��[�.�L����P��&�%���%�m�)�0�1q���Q��j��,�݁#��]26~������;	+�qE"�^�*�T���$?)@��dK�Ar���P����r@�Z��Aa�%)c8�Q������t,7/���Nx9�'b
T�e鷍��!Y�B%�C4�f��-aH%�6&X�W��:.�n��dㆺ���k�W�2��0����ͯ]x���$V<������nE��gS��4@���P�è�̰�qʗ���g�YEF<��#	}��%��S�{��-(IHt�`�������/䇎�k�6^m�[����Q^h�s;a���c�*���/�?��{	�=y�^�y}�
����?T}�U�Տ��D>��ʠ��8�����(�$f���������n���`U����<��.�HbpT�4��M�K�i��L���,�z�@z��{e��R�G�d�vG��j�u7U���N}�e���#/Ĳ�1dV��ǲm��[G�²�������\T�Lބ�w��i��Ҹ���3X�ت��i2n�D���,_�"R�'��<��d_]Y��R���iv�Y5x���I��l`�|}����#�9��Fjz4 '[�����(0م��Xq�@[�O�<(���n�@�C���{�㠸��ؒ�ؗ�r����/�O	���c�O��JU�E��.>ɺ$�+�!'�1仟b7^[��;������j����� �m.���-|)���f	�}��㮐����CE�nq�s����X����^�m/e�,��o1Y�=}LX>�4{+���zvf�`x�F�:�6ߞ�7���Jr�Y|t���|�B�tO��_��r�2���إl������{pz�*CVf[�Rb1�|����c��ю���sc_�!m���U���e�W@���ߨ�a�i^<���OP�'��h>Y�_y�1m��V���_��.�KÏ�Mұ>�*2r�g�S]�](�<$úm%����o�t9��gڬ�����y�G�έն6t2 �4:pN|b$�Y�&��U�ς�V;���]���fh�b�����xUD�!����~r��a�*��Y@_�^ӭґ���Eg�@��97pØn������&4+Ff[D5�=��f�/���mC9���r?�F�q�WN�� �K]��J��J�aw��8�+;-s'��t	�ؑ�6����$�:�uv���3�w�mg���	���	��,w�v��H2�9��v�Ő��s��ߧL�I�|��2۠DJ�8�E$ԷPĂ����bg�t��zJ��
�xE\���Z� K��S;s�q�)��{���=�=������Q��
Ƶ� ����>DE�j�GŤ�< �l�wޥ�=�:�s~��6�k��?�aj��G�����G.�&�]�O�,��w���~Mš��7\��Sm�h���E}(�-��|��}nמPZ%M%���&���^_��G���.2*�<�'1z��� �&�e�_omv������;U��y�����~8FBD6��z�е�C��I��W�0p�M�P�,��h��d�"�p%H�Q[@b{��`�׾X���/a���a�̋+�,4�64Ȇ"�B�.�ԑ��luc	JB{�b2�k�N���F�	i��CJ?c��@��c�~�k�����E��A��m{�3,��]��
�b���s��Ws��=�=��9ܢI9���x.X�vjP����חN��Ǎ�\s��a�s��Ǥ�����*�y�*�A�d\�y�NO�>�m؄DyZ����=1_����c�z��a�O\i����t���\�N�2<6� �M�����R��]����<���k:T%ڀP��-����MF��#�|f,z�Ւ�+�3Rh/�2g���W@�\oI�O�H��ө1|��v�Dd"dS���1$���^�4!ŋ1���:nB�X.�FB��E
�Ǹ4d��n�3��o��C�?��j���Ĵ�s�QPu8��O:TD�K��Ǔ�']59�q\��1��%%^�=�ص�h%��g;g�D��bѻ�V�.%s�F;L4��,:��������:�m(�L�k�����{~�M���NkaF:��W�r;$f����W,�,}RJ��_���%�+�!�����$�����%�%��>�ʃ�t/$t�����Ě:ek����|~
�nL�A��@�؝�`{bx��eD�8������(ҭ��{�p�QLbڞ���u���SXܭ2�'q�+�7��+����M�"��k��������s��*���j��A��\��cו͞&�+N��j���}S����t��}֙��Ƨ��F8Z�H��YG��k�S��W���$��m����@V�ZE�w�2��4�������_�|gu�Hɰ�{7��^Fl�����q>+C�̪4kdР�iC�047��$��c�;�|���C�A��"�<���&�_e�y��>�_qt;^Fk�a5�#D)ܥU�yl5b�y���Ɂ_��0�Ҕ�����-�������c�g��������X8 �(���=j��yȅV��]�Uw޻��.L<�q��I�E�K�����"#ى�	![&m2:ŷo�����a��-�<I��;�թ��b��q��(M�-���l�t����rBJ�^� ���M�oƖ�C�G���U�����M�iBx���`^��ŷ�%jL �9��F���T��ln�2nn@����4�~��t��z�;����~���r`����C[�uU�z�ӎ�����2�B!h^�3�v=A�>��Wb$���FVY`����(5Ѹ�G�(wU&roQ_�9k2�0��=�a���H����-_���׻ĩu����K��i�u�r}�v:�{*��|��5 �"<�T߱�Č���w�n�0����a,���\�y�c�aҾ~ߛ�x��Z�������$�����l�<{��	$�n[�6 ��4�;U��+��������G�Zr�Ul���A�U]���Q&�J�:���?l��V�WέZ���|7c��'� �b�$s#���O���U�]�Ǜc�zyi=m,���e{�Xf��+.G4J}�<j�fl8S����F�� Yv1kP
��؞��'�Ο w����0DS����wmȓ�փ�0vRM�k��@���Y3��c~�*�ŋ�~�i�>�^�x8I���W+8���.L��뮍Ǯ!���+ť&&#�C�#�[6餟�2����<�'޸e�h?äW츻��&�����{�^T\I�#���"g����~�*�^�S�-,��᭧ɾ[ d�NX�'WI0�a��V����`��kKH�T`,S��]��1��-���Q��O��N����6�5��t�¦Del�9a7E��l�O�1b�O�h�CS��sx�Ë,�鳑���s�lKvu�Gp��;(����mo���+^�̀*��Z��r�Tñ6GX��dQ9�-���@
Ƽ�����V�����;�5rL�'������;t���&Y}�>L$łp;�<�.�m�� ҭVR�����P0	�䝜�@P%���0X�f$�`�w���.�%�%.#��hII	29�1&��PjR����	.����x(c�jv�Z�-��§�$g�Ӑc����Z�iz��=�u!ܻNU��H ����g�c��v�tkw>��U瑠OQ?f�<�l5wQRaF��u�Gj���;�Y%U�[�CwD�u�n�x6'C��9�1Q�3�h��K���C��j���s%iF��e�;�k^�.���mʥ�Ϋ���<i�n{������զ�+�a�V�J��6����c?Ux���$�j�o�vj��6¸b�v��m���:�C��-b�I������V�8��`'M�|7���Uc�Q�x���+�����Yҭ�tmh�c�(�#��_���s��7�U+R�0��[���I���Ab���V�$�L��'���bU��z��Z���}HF��m��ܚG�.�C��u��UI�?�R���_�;���E� J�p��&a����X�*�"�(`שg2Y^�����Ȉ��op1�:ȩ�H�D�5������	f؅�N�m�dn�;���a{ѫ��A���]*g�]��Fg �q��J���XT`��k�a�11W}��������$#=0���CH�\�*���@EGO�ˢ�`<�������Ua�K���R"e���e�HZ�Y�q[�������+Ցs���r�H�>�_�FP�LV�9P���YRPr�~%�D�J!Ԋv����d����75����9��m+�̥[)aX7�цdDH���:��aIU�@�R��������3�9EUL�!� [��tE5����P��ʔ�,$��W,�P�����G�����˅��!��MTJr*WO~p�4��ܲe�@�oNci^_:Ÿ*a^�J�x� u�.�Fg>��l�opF�k����M([��~���P`bp��8����P3{�}@LQ�K�P��o�<=�Rf�� ,���� �f6TV�B��e�?�7O�_9˽v�Y*>d�aA$�� pf#�Ry�D�?5/�����9�`�*)F��с׿'s^vmL$r��$�����gy���)?H�=��p�_�Y�) �}�}H`��GMRC����[T���)��Ӻ	3�
�8۷$c�Sٯ4ŭ�v�
 ��	[أ������O�*}���s�S�װ����	������+�J-�D�ƫ#�SYQ�T���zBR�۳�ͣt}��(m�2;�P�k�dT|y
ֵ
�����N�
m	�P��b�tWdӌ�|$E��w4O������iUWξ��%>7�D<����~o�$�շF�	�w�b�u�R!��~�0���s��L3+���%RI�ʽ6&�o�L`�XQ��EzC���V=�E8�hu,/~3zB�.���\�O���C��5=�u�|�	�$�Z��_A��@�)qr��Y�,�O|���§[���ҹ��X���Z5uXS"����J�LV�1�d>�0%I��nW���Mj5XC�b���Ւ4:��\�Y�pp��1)-U�/�7dyE�`�}&{�Mŀ��db��\�~:��lR!o���tεŁb��<���Ϣ}S�+ҍ��ڜ
�$S݌���S~Ƣ96��c:�&-#~�T/.m63v/r�rgXw��� Ra�"�"D��J�����C������A�����HFf�
]Ɲ3.~F�P�?~�? 6����z���C�Z��SC}uq��+p��|�K<���/����:0M8�)�͏k�~�|Z�$���I
�kL�	�.�26�[{��v������B(�Q_M� ��'p#�U�6Zm)kOM����7��n��i#�a>���ڌJ�J.�#���Y���P	��=������m���{�8T
���VB���ט�(~B*>lB����4緯��c���_����c��^0/�JJ�}���k���(3?9m��f	�4��j���n��h<��E�&fV!5�B"a��|��'�!v.��֯$�0?�� �v�����S�?0s�}�H],ww, w������{�1L�RE`��GW�Ew'���l��P�Ň�ק2�SZ�T.E�z�V��	�_T�vG������iO۳QOx�&�,@�������ܴ)��-Z�ں��D˟�w���͈���$|>r�(�.�m��J��
�$�d�����45�Ȓ�N�Z%vi��9���b0�5��ʦUe�o�>Q�f��~���J"���kQY�X��]�F����@����25
��v%��3�LpF(�Iӹ'0�}!�/`��^�Q��|P��Fi6rE!"��n���X��_0Eg�g��\߶����#$����hl�Z���2C���	�̟ �{����`m6 jG����hR��~��^k����Nj"�(�|]tH�_�yU!�����|8`i�)��SI�S)�E�6������Ȟ{a�J![P���Q�� �&����g��S+���P��D*��C�U�o�c�"�ܭ�@D���s�jNB�N�sbre��3�wgn�J0�Ю�C�w�s[I��ڽ�)����)sF���%�ȴ�QO��rj/k�l1��Sd�D�Ni������R��İ�,�.��]GI�¬#wm���ݮ��)ڣ���7�����(_1����Y�i�e����h i۝�$}&��1styK�Y���ʂ�Gf%��(��{b���h��`���ۦ����K�P�!��~���zT��bD�U�l!F�2�ݗ�T��Ӎ�h�I~7g�7) �M�׏k��g�I�X�2��a��ͯ�j���:ۻH�����_�o��~������JA���s��n��un>Q������y��	��t���Ԯ\����m�G�F��V�����\��IE$(�ɹ�\'>3������_iOo�Ŭ'2�o�U5@�=l�g����E>���=��l9�^�K#��\ڑ��B�Lڏb�F��'���X5�WѾ��uƖ�>�a�iz�hv�|Ƒ��]I�M��և5*�;�,	��W>���`������Nk F�'z��
�BT�Q՗XPg]�*�H�,8������Z��� �>��K�y��8U/��D]-�=�zl��D�^�x��I�yc�+���=�]x$V��������7bb��``z��7�������ގ6�;����x{�hP��4��+�X�賕��IΨ�L?���ք��n�D��_�y���F�C�o��]�Q���Ctש=M]꫞2.�^�]4�9����{�jx��	*�]��iG�J�SELʹb:I��3�H�o�LM��G������<,�Λ�9"�4|y�L{՝�3Ć��6�'&�K�?�M�/��н�����W�4֦�Ɛ��K�})�E{�%D�=�q ������O؀l�!�NSi�����I�q)�s_gx��,ݑ��a�I��Y�"�U�9<������m���4��k;[�),�n�o}�ؖ&�9��?c1w1���x��i��y��B$�0Py'�7?�Z��G�"�q������;�^ 0'T��%��h\ϭ��T���k�0
����ڍ�~���{Ww�JU��ծ��+.��I�J'���N���a?�߅�+��OH�a�ߣ� 4pǳ�L����V��FS��S
�5��k�i�7���_aF�d�)w���ms k���15��O�%ԛ�~ؗ�l���Hb�=�"��ؗ���\�X6�?��:������G��T02�Q�u,ݯ�Vg4��j����n w�ᅓ��鸜������Y��0�d(ޏn�M��eP�FO�| 7���Q�Zc?,a��;��zF��=n��^7 �BQ���z�<�22��+腪O3��Kg<�O�����_�/�@&�9O^t��-�/�� $�fI��=Pi���d��˨6
� ���ٓ[
.J�n\Kv�R��^k��J1�X��Դ����#�m��h�V�<�^�_�`w�Bj��M �OBl�{@�lw��xZ��=���4�=\�#�C���f�'i�	��N�ORg�"�e��h��t�-��<�n���(kx��	C�^˙gD�G�:�`ů��b��j�V����8���:�D���1>���&��n�Lʧ.�K�Ǭ(��}��ms��]ePNr>o����2��4T6C��1���&�m?%�[H���n�C�cƓ"a��5�1p��D�S�N���A]]��b�+/▣n�{���������jz=у�ˑ��ހ�e�����>���X����g"X�'�V��,���wL!�4�%9�B<E%�x�*�b�ރ��`�9������[Ӽ6؞�<��D_�R!�Xk�-h�<��J�RaY��;�捅x4L�ꏽ�q�:�3j���y���a�����*瑻�"��׶(W������d��h�����*\�қ C����߆�=@Þ:
QH6��m�麘0��
��95W4*@l�1ݷuW�]D���DT��]�,��A���>G�a�<�V�u76iN���҅��L�&���./v���گy�p�"����	�)h/6����'܇�W�R��y��ˢa��
3��Љ(��%`Ic`�:I����N��i�k��շ��/�kgFdz"�wX)9=̤�r���v��7�U�����rj�t�^�;.#�~E�a܍Z+��{L.`�H��v05���eI1&7�=�	�Y0��g~���Gm֎w�3����;��Ul8;Sk������/��iͩ���n��c֙F�G���+������j͆{Mo�D� ��i�l)ɺ�)-=�1
��9rE�2z)-l�Y��i��\e�+��LO|Hs�?��]��Bq i��3�����~H�ζ9Z�8X�q�|5Jk���
����'��b�<
��j^JeՖ�`lh���F�+Іq?n)�_ۦ2�:m��?��� ��K�ƿ�eE%�o޷�8Y���+'�ƶ��X�I�@�vE4<���bWR@rC��^��=~|񦺬�Z`�Md�%���\�Fb���>��(�:(*�I�m���c�!���2E��t9����"��D�QHQ�y��zl� CLGEn�����S]Ք"@EN.Gt���̇�D~�[��p�V 2D<����o[�w�V����#1�3m�m�)%%0>@�f��BE0C���{kv���]�4iFG � _�/�@k��/�ڙ����f�-ధ�烷@P:4X��єLR/��\QO9d�D�8p�˪�)m���p�O���.����3cH@:�:C/��>�l�؋��h��9�hȴB���>�`���h�G�Y�N�ţ�	��4�	�;��ƅDҮ��
�z{�4���ꇣ�pWӖs���!X��U�T���Ԥ��z�5��g(
��J�R��/\��_k�Z�+�򂸽�rj��%,�r#&/����5�p���E�'����n��_������H.G�ՎQ������b�=Bۋ��K�E)�� ��:���@����ش'�b��p`�o��.�[5c��~&[���������$j�]��ix��wY)�Ǩ�ޅ����0����0����E+��ޡU�������Y/�#�*aB����2n��o�.�����:E��U�����:�'�?߹�����M}��#j�A_����'��يB3E����5��<'z�g�]��ɠH@���T��*&�0�ڴ�#�蔮|�̴����Ćl�Pe�2��"�c�3w�:���q� �y��|J���;
��@)��?�OO���Ao��T(��(k��l#/�����
UV$�^��6�ꊱ��$K�Y~+`?˲-��Qu�ۨT��+ug��E�=~I�����*N��r/���3~<+)Zˁb�U�K�����rV�01��Yhh�E?k�����w�I
Nm�n;�e@��J,�2g�����k�{��5m
��N�}����7�|��[N>�b�"úҖ��A��uHvGS�drW
��5	n�D�;w�B�:���S��S�s�;��S�/!�����G��f+5쐪���S�s�L�:-���P��0n�9wN�<�yz@=�c��1a�6�J��f<s����E���ӌ���mX�ä΄�lM����;�;�
c���w;ZqE��z�Ytpb��|�����.g?�O�3�b
�e �!J8����2#0&�\����$\�̰YT1mO'����"/�>si�g"�ɀQ�	I]l1$�����9|R,�$t����C$����t)*a}0D��oV;2�*�s� + ��i8��9��5�ce�i���D籅��EƵ.�����_=/��k{�LM����CR���Ę�X>+`W���o��۵�l��2�0����`�1��ߖ@:g)s���W�;dۙ�8����H-����W�'����s�sB��b*����\��m���D�C�\�|uV��RE7 %� ��Ga��\#����S�Mlvaŵ�E�b��i�������P}����;P^]���~���p�"��(�q�Jk(�O�k�	e�B4��UZ���]�L�s�'<��~`q)gC?�1�G���`������%̬ �$v̬����m��v�D>r�vm�-ڀ'\�-� ��_��-��X���c0�ǎO�@�Y�K>�AXL�� �����a��LI�w��)ع��/ų�g˹'�0��s��w�,ca�d�B!Rq>�Q8�w^oW'�f�H���jS���hMX)����cQ�\�/��x�'���R�?��垊�F�����r�4:E3�zNj��;��%�n~w[�h�5�S����Z&�"�r0hm>����:��r��a�UW�!ρ���_Q
�b��6{э7DW��Ԓ!�L���آ�����&@A�Pbxɕy�<��[m8p3� %V���W#�q�;BuB0�}m�	6:�^���^��W�Z
�o�f	n��^c�u���G����-aӉ뺌.�;���� �@$��?����
�#��f���������߹�]��VPL,p���������%Q�&d���S~9��pBzO��� ����Ih�2O��dS�6�'֠�I�3��35F��R3����9.�#��>���ɩ��J��4es�	L��*2�3�{�	]�����j@�2f�@�l����� ���F����O0�̱��ۏ��(���)Sz@�s���q_;N��� ����Π��C�_MU�F��Nz����x����e�l8���c��Ր�Mkw�CT٧��n� �Fc�f�7M��%������|jX�G�v�17��I��&��䃿cO�kO;~$+����0��-f�B.���������S�Tw��"�;�k���Ǥ�d�����(�X���HC�c`X�^�)t2��QHR �~����־n�2���g΋&�%�����w1����
+'%)�ݷ���pKO�����Q�3� �P��@�]/����Y���o�o��l��H�'0$h�S>e�����C��ԗ�]���)��[�y�BaE�͂�_v���5����ggҺ\�m��z�VR�8Ж�n����kn �!��\�`�y�N*Uh���1�5r��0���P���p�t�����3��g���7�q�l�� d�\겛��3R�4�'c��6^u�*��SCO�����e�C���hrA�m1��vP}�Q�KY�55��>���s��ѱ|��.B4�������D0�z�H�&w���]q���5��9�_@�n����P��V�;_G E��d�Ř�<�O~���ejV킇36<��F>i �l��o\�K����j ��>ru�<�iA��s�J��bȞ=�Z׌�{�tt�8v����xޅu�MT�B/^Ej���CJ���/���naiB�����!f��y��<9z�ج��*8��u�\�j���V���B��s1dW�Ϗ,6��]SH��;Q_fT��d� ��8��ц�ȍ�$T��?�P)��6���tݓ��?9�v����.W4[4�ɟa��d[^�÷WXԈ	���n�X��|��
y�>8�\�m7���t��dֳ �a.H�8>��Û�y�m��܀�$�c�9{Pj�H�2�Z
s!eG¹Jk��L���=�$A�����P�9��'墸ۇJ6���b�)jL��؅S���e�"���Xɂ��Ɂp��.ÿs�u�8����_'-�M�О+�,��GS@��'�&/n��PW�Z�d��s��Y��F���٠ ����-e��B,+��w)C�N�j:�r�{>�8�%�{��U3�n7o'��dN4rx�aU1G�T���TSU��t5����jnHXf�i�p���l����&��Fͻ�UpK.��k`�+�vT9F�ܤ���غ��
�=�l򄹍���-C�x��s�"/�Y��5�+:�"Ћ)����ED�҃Q�!��#��׳���e��oK�]��BWm��#�WJ�5���Xn �kG��+�����<��#=. q�0qN�c�
����y���;_�@l8`��#�?r�!Z�{���]eH9�cx��Cm��d�4?ق�SF��@�hƥ^�K܍Ӓ̞E�!�l\U-���9� �Csw�hŨ���7�֕�s�f�^(te��Q�>��n�pF�ʝ����1�ܒ�Cq'��DHIZ-	j���_�p4��;�b��D���.�����"��:Il�}��o�^G7�2^�����W����鳀/p0���+<%c]��;0:܌�BC�l���k�r�xL{�������da�h�E�ћEMN�hn��=�L$���D_�l��w��r���5k�I2F�{�1 ��VL�}`h���󿤿�5�_O�T �F��x݃	�uZ�!��ĳ�Wd@�����۫���S't�5,�^�B>S�ɻ��6��8?,8��P��Jn�WECp�D�*���o������@8�E��.?�R��̶�XEÉW�C9I�a��a���=�VBO.o+YQ�7��ۃ����Y٩m)��[9^�`8�Ĝ��Rk$���Ġ�C������В��}K��/o�y8�n�'���Zu,ť�N���õ�q�Ez����!M��Л��-%�>p��D̆&=��<V�)�<C�"�ߨ*K-S6��6�{A� �,u�Df�Iم���/R�&Lke�j]˾�r�\<��ޫ|k�����t5�-BE�����o�4�� �W��Ts�^M�"�n~�L̳G�]d�����L�Q���ak��������F��´d�%���P_�F���_�1߽/'�t]�{�1){n�W�S�����<��w�F-� ܍��ܰ�U����^��Ӣ�>l�/���H��Rh�s��=�S�D��9��f����q� JY��\��@���|�\^u#K�I&��zr2�Q*��>���ۘ�=��_�O��:�k����&&+��LuB/=�tמ k]�9v�sxٞq؂sb��I�M֔O���F�B��0�<M��@����kcd�Oa��E_�� ��%w#��s��eI�۷�i"8a���)F��[�\�X�T��������R��9�V`�v��l���KH�d�U����{U��hN�	&�>���=Уr�f������s5���Nyɨ�D�@�9M�v�IEb�Hg��=���K0����@��4�l�9e�KW�X �f����~5��$�`r��m��[���b�Νl7;X�ʸ�8���м�i����p�ݐ0������h���Ʒa#����U��u-��] �O��:sC�m�'�"���:X!
j��Ba��E�h;�8fY�W��.�9fP�`�/�H���>�<��=u`l�,y�&&N�ҮT`;͓�,��p����G��T=E$�|�TXk7������R�Vt��˴5$�z��Q�y��	��aP��z�ԣ=��r��A,.Z�AxY�.]c�8��:l���IW;���|���@�V�ݼ�� g��a9P��|���I�G}�/,]��߶�Ӭ�`����z�)�b�)�Ƀ%�~X�_�����l�������bIE.z���ۂs��MB��k䑚K*�R��\}�0l&X�̖�y�=�2,��o_�cn�Z{��#VM��E���fK�z|�<�a���*9H������pBaaD��bld�?Y��(6��ˢ���,���8����������k���PP��ҍ��G��̃Jl�$�Gַ!����Y$}[��62��c��m�ִ�}��ቴ�^��۽�n����� ڞ��NR�����Q<=̏0qռ���:C��v�,@p9�e�׼�5%qf�g��ʇ.L�ɳ>���@���0N�Av�Hgv/��hˠl~���,�sH����[�۬t}U�>�KpLTr��U4��>��k�����Č���<M�0�����H�%�_UPZ�,dH&�л���P���8�~�2��!T@PV'���M4쬍���k���j7�`��ƶ�Bm0�f���#�q�q��������L�@�u�e��^���L����4����O�����+۾�������N|�;l�x�����$��*�D4Ӝ��G�7O�LP��o;�>��'�K�Gж��z�~#TUUti"Htb��:�F�
S����C@�,2��v�`��Ӈ�:��Ȯ��(W�N훜��d�854T]w����3��JРЅ���W�'�b����)g�>)Nb�{��h��J�r
�1!h���3ǟ�<fl�����t�JI_�)s�\��h!פ@!%E�T�]�-��w����iP�q�ʡ&��F,��pB���*�9iq�|W���@q��H��߸=�~M�5���o��堑����S7~`��_'¡i��4=�r|t��п��(�</�,K�H�i�ftK=�D^���tp<XR�`>�Mp�����Z=�}���o90a�{�l˧��x�s��Ͷe+^s�O�m��{�)OGs�.�ΰ�W;i�)�p�M���I�ir�AH稬���)j>�)���Ӂ�#��Y����xE���Q��0�Ӓg�>���J<�#��;�B�������V�A#�/w�z��Ճt����,�~��O��������c��u�y)Z`I*�`h<	���#U:p��j3%0ڶ5����mL(O|}�4I2�?
��V�/�T��+-S�DU����|K)�⚂��X���:�A�?�퀘o��Z}�$"�2"dc�H=�m�������ro�D���FahԌ��#)@��/7iI+��Q�=&�w!!���>�i��ٜ T�LO%����
�Y����P,2nhl $��1��{|�p���kLL���H�G �t�/�\�s�uWs����.ۇ�4Z�y>	<
7A8f�7��.L�&�C���8�*�O�����_���+%�O�1��0���#'n�Cu"y����K=I��ɼZ�c�)��NU�����u�+8�_�@ĉة�$A.���|�d[��L�c^�q68@.���>�ta#��o�+E~#��(Mm���0g�ܝ #%�}bH���T��Ak:?��==|R��S�?�������S��Ћ	�Y
���-���/�e�J��Z�K(���L�};E�pg[���,���C��̸IFa���ňQ*���!o0�$r�@��p�h����������l���k%w����𱲈z�E�������v!����~$_��ʫ4	X���z�/R��Q�w!��m���@���f/�������;-�;���.�[3ᦗsd�wnr���%���1��]U�9�]���F|�l�1^[���&��ag9/<݁I4�_}p�dw��ML�Im!���봩�w��+Xs��7۩���Kx�%����r�p ���*۞Ք��� ��amc�\����v��^.�rA�H�`�~1��6,%f�}��L���JϨ)V���.Nf�E�|޷W��Zd��ݯk�#���ND]�������u�-����&\����N5kH����J�W�"G�@1���C�b,���
$��	���A����5����_�� ��gwh�â�v��P§����}q��>�{�	Pw�F�r� 0��]�H�����9h]�Gw&Z�(\�F�(�&�q�bڟ7��b�H?�<m+����+i,��p^�!����(dj��*)�r��F�5���1#���(�6���N��u��,����FvR'ӧu;�:�����+�f(c��1�ֹ ��|#Npeh;��\}7V�$}��F��<�ȕ#T�P������4��"3�H�`&�#�W��-�x�	��	pz$��7XyYBzE6N�㈛����6�\o8��Ti����r�8K�$z��7v�	݂�Mް[����{)��Ń>J��߂����oPK�ȈҘ�M�-8����5�\�/�C��'��y�ݰY@`?g�ا�(�����c�������F﹃Nm%K-������<OQ��(|e򕋜�|iЍs��&^�H�X�&�����92������B��"�/xZwk1*��1��9��{���j
�7+݊K��߲��y���x�~����-6�E�����=�A\A�/�n=L�� 
��CKx밀�F��I]��O��)�܃A��0\���c�0^oVG���K ЁD�V�J�Z1�5�����I��0�o]x�ZmxUWx�����Q���^Ϗ"�)fO�Ja/��7Ԉ�^���0�` ��|w���u�?�S�N�JpD^F�&�JJ�c��΀
$��*����� a�m�I��[[���k�Ӧ�8�6���o�?.+u�5br��¦O�E���vrx��,��@��眤�����O�61rq?֯���[�a��P�U�~�10�/�{���ä

��.�H'Q���'³Ҩ֧4Q��ő���ǭ�i��|	�h0�G��I�G�W�?L���j�Q5^V��>ި�
����պ��)��I�}�hOZ�dCq���T����6�g��S���X��OUg9A7�{��sR��U�C@�
)��[�֩�I��6��?�96�H���*#�Gd�Ɯ��Jq��?hX�C�U��峖W�B�u�/_�
}Y``2j�w��Yq�W�N`���}�����Y�f�ܟC���`�Mw���V�Z��>�l�8�ɶ�ǎұ:Z�y�@H�����p^&�J���֐����1��N��b$�����ڈ�Sv�7�Mǀ��.0��ٓ�_�I�������pmO���2?u�����l�zl4,'4����j:g��U/aI����ɾr_�	m)�	������f�,j����W��^�IK������P����&v�,��M]L���d�s��'����o�Kl�rȨ[����	���0XE�4�����S��1r�����V��~v]?!��@_�%ˆ��s�
��,&\���4��֎���d�u��P0І�����|�I~�{�Y&]G�}��Z�7�Р������Vf�[~qb'V6�W�z��5v��Q^`.�Gh�������+d��$jJ쪍��P����¡�,"7�HY�ѶdY�-Ѽ��LM0�I�R�4FP"
.��Ϫ�'M�f�o:�+��]�n�l]�Ť)./t�;qUR�hD�wh��c2���㼼] �}�������p� �z��/�L6u�3N�|��Tl�F_�	�uFD�D�p��M�I�kRvQ-�2��y��`_���5�`=R	��t��@�h~z�Λ}�~�3�y��I����l��[����2�ݜ��):�1,��]����el厡��`y!u�'����Ew|?���ۺ���T�̯�����8��m�f�~��FR�_�0v��cxh{��q����a�~n}�i<�� ��ڊǼ��謌�>o�
i������-s�����{����Fv�v[�s2k�����j���\E�YD���X*��p�G��@B�wUM��n\�(:��̵��(���~���Ō����ص
T���	qT���x%���6��$Z]���e�>�����r���{���^THd�]��XN��	h��Ql�;V�&(mZh3JP�>i�Q�<����rjY	1�ʱ"���pQ�&��|NҖ�k�����x�2w��s������X�����59��:!$�_7��EWwny!�����ĹS�����y���j}0��5���
тũ�\��:-y�a�H��K8�@��`s��a���`�ʏ{V�[5�����P}7B$�깊��}}�4<��|���W�s�=}*}�mv)������P��m�0�E��x�L��'К�p���Ιm��tx`=)�&S�8��$f�^����IJ�c��3z�&���o�f��=���Cm|1Q��4�9��OA�v���$,!�<�:C���?^�:^D����XJ=-?��_&q���'��C��,���]�4��� ��g�8�'3s^L4�gk�(����Z5x6��?d��4�G����n�C�O�>h9�����Ȁ+ �񊺊������[Z��s<�u�2�|*�z�)�!%2p�Ml�N{�/��݌������HaA�,' YB:d,@��(�z|�/C�g�s�` |��z���SXO�믠5�F���,���-�����0P������$:���g��7 ;=��G(,5�d��!y��xZ/*��	2��/�竁�[89+!0n:���W�r0��_�bns���w�-�k0��WF	QBۍ>��p-Q��zm`�KO[Nl�r�ɱ#�H*�mR�q�P1�D	�P��@~�y���4�.�aD� \"�F���lJ�̈�;�⠤�"6�=��5���ĭ�J��G�8���F��+?�,.vW��x=r����f�q>j���\r �0xD6G�;qw_�H����B � (��|���'�<8����o#��T����<?S�8��p q�Q8'r�9�`�S��i-Vx��x^�c��KO],���>�"��s;r�TnmG3�v�F>z4�4.޿�Ե�G���U��N�T1VX����ʃ�18CŒ�d�>�,0%��v��� �b��v^��<�D�a��A��2��RoH�H�&�U���2���e�-��s�����{�,Z����i�?k�9A�y�aӋ����/h����3��0�'%C��&����"������xJ/��y�To�BI��4���;�+B%��usC_j���A$F���|&QFx�������ȶ�������5�7���	��<%c�M��������a�<^�k�;n�ߪh5{<�����a~/OJ��f�g��y`äe�w���t�����GZk�l���<	�翷X(� ���QmÏ��|��Zi/"_䱂��� �������H������T�m͘�����S�_��K��N�;qf��n�����iF��m!3�,`����C u���X��4�G���E���ۖ4Z�x�,l�N�/i��p�4�F���K��pZ}م�;{aY"L�^������E�ˍ�����}R;ªe�)'y�b�/��	��9���I��>�U}frR0��,�
~���Y殹'������f�*vc5�y+��S)�r�u���z2�dQk}�)W�G�ZޗY��0Џ��K&�\�@�Q�Î�	��Q��D��1TYOn�6��쀺Yh��R�$$u��i��Yx���-i)�u�: ��֧�>�PwVƯI��q����p~������&���wj�Z��,�e��@���_е�G�T�O���qiɺ��}��UpGʆ�	����6Y�8��Y�⊿�N��Pj�^��j^��zW,Q�C4K�#~u�C�Ԕ%ó��&����l)�C~08P�R�y��\��o���ޜ�EDC�4���!O�¿����҇��ߨZ���ۑ�܁
˄�UU�}��;ٛ_�+�i�|8��i)]�����2U��3�g�`�v�l83�[������\�������Bo|�~�v��L�-����Su���R'P�-�+8���Ǥ��[B�~�>�G��$���S��F����B��iq�lozհ��Hx�=�`IK�Q@@*�p�P/2N�@�H��rZV�]͗A���3���p��.��\�ף� �D��y<���Q�"x�<�J.��l��T�K���:�S���`9<s��9x���_��V�P(�J�LH�T��,�dL�ͣ�ؠ�tE��z�ym�PS�@��p8�Ev�
����k�7k0��7�K����Si���VיB!�m��J�%�Q�̓Z����Эnᮚp�?���{@�G��Ҭ~��ӤGR]��)dvhwx]��Ƀ0}�KSH��u:;2�$��ѷ�M�5b7��5��s�n�?��,2�s}�t����ES�}�f�G�mш[:����� �[��L?��&��Q�$>'0��ye�J��*�E+��J��~�l6�UhAb^� ���Ņ!� ��!��'�nSJFVa��F4�	Au�:21己Q<�{x�X���5�B�K�a�H�1bM|a�zy�aǠ����p�,�t�op�	R��������(v+�}���\ߕ�a�f5̑�p<���"����-�9�fw<��\�go�V2���� ��1�D,�݅��Ǵ>�?�Y˘��\\���>���塯��|b��ܲ��<�6rG���P�û��P<sj,��spB��݄g�A+�Hm�\^�9#e�o�nU}�k��c�E����,�Oo��u}NG�!�g\�������$���U���P����WȊ���Ip�c��~A�z3g��ۋ. H��{��!GV���zT)��J{��=V=��Z�R����%Z���i�����Y�"�kZ�
�d�U���$�ؼ��B��=-}@<e%�:2�;MRBd��� B�
��c!)��PU���+�=�xM���iCu$��Wj��[��z�LT	�si��?G?�K/�����sUcc��Im�ʽS������$TB��xOt��5F��T���)��R�W�s��ٳ�(h|�����	���KGzU������Z9�?��m��I�
���iFcyֆ�+�o��U�k�t?;��[m�]I����>o�˭��h��T�]^��"$�#��ol�`�L�^t�\<�J��*����hD�������4����軲��@@ ,B��C(�(O|3l{��t쌲P�[}qY��$"j-Ŗߚ$��N"�g�8A��5ќ5�5o�Xe�W#��;��o]A�J,<���X>�X���'��1���"B�ٖ�3އ�SyZՕ�n�����[���e��Mg�r�+���=H�z��L�����pKS��� �a�e�{����Ԑ���yV]"����ؕ	��C� ���R��O��4���)	�:%
l�}�N�
�+s��0�-���A]���]Y���i�O��X�~T]�&-�*>?Gٌ�Y'N��S�#����݁��-�աYIˁ�p��n�|#�8��\vp�E��s����{����KM��el顋���i;���$'^/4����t�ޮ�Ӌ��f�l�U�� ϛjrr������~�/����NN�:z�ӚD�Ň�I���3�Qaא@�x�h�hu�v{˛��@ }����B���i��2�Tsw��U�p�mU�v޵����G�q7��ճ�N�5��g/A#W��� d_��0���!�>���*Z~�4������P�}R~G�+Ok�U���}��Dv�rb�a���-J�n�Eի�D�H=�6�5��L%�<����7a��{�X�_t�O �gZ���.�/�ړ��g���H��QO�%`��DqQA+���=@M�w��";�r�}V�7�k	l�d������s��.?.X��b��k�ע�j~F�'p�4P�o�[�� m$d_���J���TSt����/��7�ߙN
���t��DRv?+NU����6���A��#���D:��Wޯǖxiz�UK�����g�=��)��{c�3DX|��1�f~<����.ў��*�Mwm&g��ǸJ�O/�����-]"��>^l�1�<�v�D4�/'����r��|�,܋C_��DW�[X-6|��,�ic�$�a	��ch����9�\�wb�n�pY��3	4V}Š�O��?�a����9��n�Q�x!�ŉ$H�xL����7�>������᭔md�C�pI��ƅUh�g�IV\Pz�i�Y������3���G�� D��-jy�c)���ۨ�=� @�q A1EG���|�j��/3�U��e�Kɗހ��n-��EԺG�Y�-��Nn��Ʀ�F��[��E�Û��!Zt7��DG���\j���m��T�Q�J� �-�e�D�N�:eh�k׏ B:56�N�n��<�����$}�F���O�}��N�(�DvT3)�mRvo���R����4XV�{a��v�8�$��i�1�r�yc�~Y̧��9�[����z�bm}X���P�7����'�B����۬l?.7>��@�W1�B3�M��ޖ\'&��U�߬�6�<�IXsn��4|�D0+�����/?E�	x��?��FtM����3�Z�
�m�H�����W/�UH6U5,
q9>�L)r�b�R��y<�*����w{wՇ�Y���h>��ѡ�/���s�MtB$��>�Lz����z�� �I���K\�f%C)�s6� T;�
 q�iW8".xh����i��$�M5�L߫�s�&��s�����\~Gfɞ;	��9g@�p���"5|o1�د4Dmm���0vlE��\�����n�*m���"\�2�뵡��m���_H`N�W�Ŗ�J�z)�%�{��n�(-�J�����_�_i+���e�_-����'����f3e�Í�K��OwC,�X��?o٫"~P��h�l&�B�|)g!؁�U����ؐ8��B��lG5�0_����ߵ���곥-����×\xb�E���˹( �]����
R�Ġú��u�Z�1�4�0*ܻ�z�0�j�H#��U�]�
��n�@�ђ]<.���j�s�pÀ��T��(��mF����(�k�ʈ�
�m����)����!���?�,�mI[Ls���*���M��^[\텍��e�հ������f�")���+�c���w�]C��7��񕡜~>��E�#�:F��E�9W���/z5'�*�Yr\��41$�)���(%%/J���v@ħ��b+0;U�Pa��yD�2��LX�F@��F��h+5��K��J��@s�FVZ�8��R�`s��T!��5�o[��'q"?�0��C��i3ӂ� ��S��G�> m{K��N�(
^f[�
�vf	��LB��8����v�̌8��o��!����SHL�^_c��A����%\�S�|��V�����ꤚ�O\�Z/g�}e��3UJ2�>n�8r�؂k	�p�WmWJT�ڻ��G��9�9�<`%����D9�����<F�Q��EP��c�"��뚞B֌*\k3q�<�T�i���<s�Ji�n��%��ե���9s����m�u7%�e����q�5vO���'�x��Rϋu������>���@�������F���+����K��~�]���0\�mK���_c kI��?c�?�N)A�(K?eE"�Lđ�M&�d�&�	�=\z����
��(RA7>���� ���$�8�$�ƈU�K*GXͥ�Y�%�k۳�Q��*���x�~����$+p�����(��6����+U%�⋓�<�GJ_E�.;e�iˇb�t+%$4ɂ�
�6��t�p	����G��h����C�F���M�	���k��Q��	�_.y��'�w\��1��7=������M~����i$�v��E��� L�S�U(L� 5/�λ����K+��`���ԫ8e`|�$Bمy�ڙFOD����L0wR}	Ň��	U��r�e/&9)΢������^�,�u�@hO��O��0���%�.������3�Rg"�������TҘ���Ay�l���
�n E*;p�ȵ���]Á:��9c�����)��HT�v:�	����ɲ4O���m^�B�m2&4I���tE��.����
������݆�@����c#���T
R\2����y��
��$1�2s�
by��(W�&��Ɉ�=�U1��q���k���zM�}�E��U��:�_A�i5Yi�hI��˰��L�#��sk�罓C�ޛ� �y��1�*��7��Oh��s�ڤ��#b��~�l՟Sj��/0W�:v9}Z����Q����cuE&H��1kC��/y��:�:*.vLh�����p`Ns�h��ARH��{�=S\^3~��|��ٝ΁s �z�A�!*ܝ���%�J���1H�]��X����(��� O�fB��-_��6��$<�5~ޓ�6��V�����녱���Qx�[��OC��E��ْ�WH�d�,�Î)�O8�=D���v��3�jVU�w�'`JHp�Zu�v4g�/�(N��9��_ƚ��B=�0����'�\��c�>���7�Di�r�#5�"K@$]/���gЪ�n�g.���<H��Z����ل3����f�Uxz�,�IMQ�U�1Dg�u_
��*)�� ����D�h'	���P��26.�u �P&_�5m��`$�I�=��q���dg��b��
��k���<�>6�6�/l{j�{�o��KJ /0<T����=�׬��i�F<�.��;!�続�4_�Y?�W�д�d�\��Jz��"�D�����'�?I�����[�_� ?�m���_$M9g(���duc G�j�п������q�:��"
l�-�w��o���������M8�]xy�=>�?[(�
S��z#��7>6�z�C9=��ω?����3�(B/A��:2���?O)�lx�n����oR����sdl�s��Tc�g���{��Mh[��՚Ꚍ�,��v�!~Hy#M�,�F�E�LS��>�^Ch��j�������"CY���S�9�Oz%�bN?���2'&��s�%�Է�����K1�P3���2u$�lI�5��I,�s?YmB��pI�C=�Kh(Ì�C&ꖥZ�Df������0$�(	o
������ ��gB���G��{a׃����%#2&�����1"���1�̈́�'����`�+�K�a��!�����
�7����d�7����0�Tb����榺a0���i����_�1U[9����x�� Z���)Ĵ����s[+\0S�v��v�I�M"�ָ����wǪq��U�V�*:B/�)8Q���1�-�o
_|S�iA;���7���J���*A��$�޴�̇;������W��𣫧�ֵ�%�#X��r0ߔ"W��	7�_����� l1]]� �[�0p��f��B�y��a ���y��_5��׳Cz��5���p���Ez�9����']A{	�M���e��b����x�]�YRMW��8�?2v�&N�����^B�̛;-�k�`Ĺ��nJw����Lt`*��7�goJ"CA����5��NW�y���rდ�H)�4eP=� �~/����gz��=�~�y{+���+嘖]����^Gt{F���,Sd{9|��=����x�i��F#����f��ey�{Ӛ�V�����N�C��f�y.����s̓v���]-/�"�\���Q��:�e��[�>Ѹg��A�Q��%���N�\K,[�r����E�o�l��zs�Nn�2�$��3�eK1�i�����
G����j+T̯`.�G@+{=c7���\��٩
~����J8'ݺ�H�(g;�8�4<��~�������쪐�5��x�Z҇�m�ڰI��m����D�g���Hutpſi)��R��<YA��\����m!(����j�.d��v.����8ѐ��q7�b���w\�w������#%���V��?5���D]7ܷ�W3���J!��&PA8�Ӽ��%�/�mT��S��s�n�&A�lw �L�#�'r�	 �jY���?)���H#bܱ��H���Mt�ޤ���=��� .��h�Ň��S����Ep������H��yJvs�pf.6�@x-�|�Y��8#���zɯ�a��G���)mJ��8B���B�b_���(���B5	t�RH.�^r�ĔQ�2��ߥY?hi�E�k!�Bىd����u�ݱH<`&b�}#�H���2NQX����ϒ���U#
��/sK�$g��UJI̚QB'f<,�2Y�<E�V}l^�Q�?)B~'��soY9���}qR��l7 �$�l�_��V&7v*���y��;��*���e)D;O3���?��������N7햯"OR��M�
�Ɍ�^���'�`'TuQ}d^/��6�� �u�ݙ��P�+��C�A�!�,**�i�@��@����{V�Ft� =����(�����9XI�(@ ��O&��N�~�o/`�_��duKÉf+N��ȭD.V�?(��[s�;:|�3=����h}��(��x���i���n�5^���Y;ܱ"𲧜?$z������s�mV�`v��6Ƕ�=��v��?�Ҽ� J�%��n�?�b�"^�����%D�������A�b��.U��ѝ�)�C��u�8�l��E�'�E+&w�;�<z�xN;>{�m�&�����3̊8��f��2��N�9�A臤��7�n��w$��"��cߨ�� 0��ǾA�*�����g��8�;b*j "uWE�|&�v�	����bg�Bj���R��SDp<�~��Í3Nly4�ߔNCgq]�ċ3�����-р%���nTCd�$t�[���{�,O�_?���wbn�����L_"T�� �(�եd��J_����g
vhG������dub��g5���O/���=�����	]L�Ƀ��_����劻ˉ!�MB��Ч��Am�j�`����gڋ��I,*�)�?!��1M|@�/�����R�7�G*wwF���QGf�ʥm���#�g�4(�5�j�<����WxU����}w���)��--S��1a���q���M�bh�J����3t]T8���59:^o�{Y�?��\���d]�T5��d�W?�f���.��֍P��a��X8����?���Z� �l��ݧ ��a�a��E�W�� ���E*��ҵ'�ʪb_&{l���q�8uys��ݑ8���0o�~k���
��r�"�Ү��aj#�#j�:[*�w�3s�[K>��{@G<ٰ���+��Ը�K,eIe6�QN�>o�4v��⿻չ�!|:A�K^�_�
��?<m&����'��$� �=�����4h�����m��G��=6�9AR

v

i�M�_�ߔT�b�����)5+�����n���H��ȃ�b���|r��L������?�˿�acBɮ(�ӵ����*g	c�.NmO^%����I&5����tf�n��7r�)�)���7���pb%���k���zMhZ�˟^#�`\S~vRhg�#p�n��y����N�B��R�#SY�-Eτ����Edx����qG�ؐʨ�ۘ��.�A׿:�V���eb-zey����Aj�����+�V����9*�_���Y���c�Ő9���#��gm"�x wqI��V���3��|�s�B�	���
J��^����D�����5�8$!�D���S=���j��7�%�b���B�r�ɞt��t��"�����U��'K�r�~��u�h�7cN�3��rLn�uw߼�n���GC��2{��Q��NT��:��fd�b,h�!������&��x�6Ѿ��wk7�*T\�N�2l��N��oٶ�����A�C�w�$<"^걱+}.ҒV��K�a�<+r@�[� �����W�8�I�o�6�(�lQ�dPo�/�ّ��&���p�G���U9��!Su�;�XK�
�KR�ư�e���KP�B�^"�A ���]��a[�?H���̀5�yX�o���,f��8�c��P���������V���m��&�Rdc�{�E;�('�n��@�ܫ�L�{�eN|ǃNF�2�-5mq��ѐ�Y�`���4���K��mw�Ӝ��	Έ�K`:;)c6ŕ�]s�>��5w�V2��C��5{�}�$b<�ZB��[�X�ࢺd��kbLzu��`m�ԨF������Y��	��W��a��2{o
�����S�ݫ��b�gr���.s<��)���F���8�����cI�[E�v�p<�Ja��0vy�J� QR�rr5$0�x��	
��^M����5�@�lB�>b�yKkE���S #-+�g�e͐�g���IPώ�/�"� ���e���≺���a��y��p|t�m�����gF@��eb���Dd2>�Kr!� �#��V���L�5�?ㄫW��<�!KtSK5��5J�[��<��f����	#��؛�f"z�}��n� �݆�ggƐ��/K�ޱN��M���P���f�l�-��u[�H5g�����vDJ�E{t�'�R�ʟ�=ΦuR��\��ɬ�&x8�X܄���
e爝���}�g�[����sC���$��0��$σ���6���v׽�$�J�7�--��c�j�Π��Uu��z�6v<~�� 5�t�9�S���}`^-das!@�`�0�^��&O՘C��
�$oѿ<�A�|tG��$�w1w����t6�d1�+�
Sa�Xb(cH.6��p(CJ��˼��A۬��+u��ka<҈�.|t��'���L; �5�a�'v�I�����Ck8�7�k �����p�����Q*�?�� ���D�>���~�' h�G:7�*�\{t��鏎��8i8T���R�VHH%�Xh�����sRE~�v���-�'��N^�:~�!�NWLޅFv�s��%��
93A��T�n:�gD�Yer0PC��v�-Hf ��@�s�4u"�t� K+m-bXu魊�Ig=h�TР��Pd���9k��=P{p��`ߖ^=N���ސ�����^��Z���^�fw�~x���6;.���E��c��+��B��g~cx9?��~bOk�;H�)����Ȓ*_��uѤ��CR�F��2�[K~�T9�-R>�T�m�f�Z1�͑���~&�V2�ƀPs(,��F%��<�������Ld�_������-Y��0<�h�k��4�u\��]T��*�y�s��Ӂ j!։�k�pu3Q�(���'�QQ�E����G�y���U�t��x1�y��J�}��o�5!e�����9�UF؜��j�ӂ�=���XE���w\"���"]g�m���L��%|���5��쳷���)�ˈd�ce5w�����i��J����[th�8�wᩢ`�]�$�2�W����&�N�]`��0~�^��a�c�H��ʈ<�?8,�nӻ�RV�9���:��UW�t]�5'T��l�g�x%r�]�H�i$|ODH���^�"�֑�U�D��I��ɴ�y�bE�D� �.2+/*����β"4PY�7N@�j>�C"���ܬ���#���
�&��0�~;̠�υ�h��G�Xh�z�
��7?H����5�v?O��&�(�Ժt������q1�W��v��q�D���?0�D�A�gVNz�:�>BY��oE����&�_�!��+�Q�����#�~c%j��[�v%�*���91���J��ޤ�D�[Xw��g� �u�&�g�R���q���4W�j/#���^vy��M1�72�@�r>E®G��S�:�D5��s�#Ŭ�y�0/�����n�k~m�����;j��83L5%�B�wd�7�^����;'^@�6Og��{/�����A�p��d`��\������$����X�Ǐ��A2V�����������R���L	g�� >�\P%��<a�$�P �ߵ}�9�=_�:��c2�{��|�A��g~Q`|V�������?����©>_�ſ��}?n\���t(�Q�&w���rîi��Yt�
�K��x�$�D���ʎfx���l=�jAc�!;��C��9��-���Wi�2�ٍH�Ú�z�J�\��E5�[�ʊZޯ��e�y�Cc<����y�����HUgN�s�bU��Ul����H�q�V��̊���e�"�e�kb�yj���lB���Wm�S���17�+�X�U�S�7�Ջ�~����8M���^JP����c�?�jП��\W����N���T���Xxc�j�R�u����<���e˽#i�S�F9�^|�=�Za�vT�|jOs����$��e��v2���l*�j�s���S�����Bp��w��ݜ�$p�h���yYL�8٘x��C�ō�,�f��3]��kۗMGa6�ވ[(T+��W��X��,��X���w�J�RR8�ei� Ů?3�Zp��~�=�>��xC�����Q20�Z�Մ���q�����ǳ"Ī�1�M�v�g͗�w<��NA���0<1��,�Y	a�x���A������P3�r��Iΰ�;K�M_(�L�p�TD�߀�&�k�M�i4V_�����ఝ�΂�Fr�����h���,&��U� XY����ig��\������5�C-4���,>t]���[�ca%�;]uـ� u��jet��h{/]�n��� g�_Jl+��)`�X�oJ�#�S�&�`X*9d�ڹg��Y#Q��F��o���K��aѴ�A�l�H�4d�Ҷ,%y��+��G�%�Q�Vۚ��N�2[����j�x�,�F
��	��|���mo�����BX��O������8�Vޜ�1�!3A�q��aE�\��w�����H����;�
�yB;���[�;;�h}g#WT���F_���tՅc�P�){}��ƿ�% ێ���EA�|�l��Y��=�#;�`3����ް�q��/�V����н��+׾$!��}sn��*f��B�WMA���G2h�'&�Ӕk0���>��F���As=]rM�i�+���K��Uof۲ �5k0�<u�i��Mp�⥗&�5���l-|ltX0;�Ȗ]���^�!�5y�h���|ڃ�V�a�Z���S���>i4����%�����F~Z��&�d+���}އ~�)��h����N�oipY�J{U�#���>wȄ���h��}._�}a�(sOC��!�����ƚ�m_��M��y�v	�;�J�'�^��{BZ�P�n�+&s���3���R�ǧ��_`F��~���9���X��\0�q��y��Qw{��o&�t9�y�m��TX.��B����2���qz�e�+����-�U8�#����O\x�Lk��E�ҷ=掹�?�X���`�ʭ~��Kֱl��>H�n��[VfK��ǵ"QV[U�d��L�ٗ�U�C�,o�t������.��zw���=��>%jÿ\�6[b�y�^@9qy����8��[R�7T�Stt�-.&,�g&�ĺJ�*;x�ۊ��M?�3����F6,�� ����?�sץj�[K��m]�̼�ۊ�#�_�b��;]�P�Ռr�Ƙ��"������&Ц����dt�	�`��R���9m 1Mu7�&_��)� >�yH�ĲO��=G��S)�<YP�uC>��8[NG�4���b���DC��Ba`�*��������]W���8�B����}��+���`5*�;A&�3�w��rλ\��`�f9������*�� ��-�V�2|v�Az�wB_�P��uw|\�v�@�ր����s:�Q��(����ɍ��U���%�Q�k]�eNx)/�%���WoT5����`����p�x(�yw�i~1q����B:u�H�&'�B��=9�Q�w�1'41�5�%���	����5��p��'od��}7���=�� �������Q��BcOr3�*�/��	7]^9$��C�7������ B��2}�4��x�du�Kɋ�u1�˳5ot���\����oZ�!����Iƒ=a�L�|��7�n(��l�=���@������Ӄ�#���7Z��D��YD�����t}"ܛ#��7"�C��#�4g]�T��������aM"���@�<\��]L�ݛ��qX[6XRj1��ݔsE{޸T3���._��c�$�y�A18�3$�&��'���dh�������V;���2��V���d;�Sf߼��V�<�/⊣���?���p|ةx�k/���ږw�$8'� Z��Z0͒�9�<{�T؋��F��xB�i�OA�������_� 
]��q�7��'���:�D��=h���Se"���2^t�T�>XqZ!�{N(��y����"Tm�]��D����x�*�<��wPX`!�9�h�ԫy2w5>�E�90ֲG�^��~�2�z�,V���o�"	rw��D%�!T[�Lҹ���������(�v�5Ԉ.�RP��:��B��h�²/V/��~�|�h�5��C���`5��ʼJ���K�b<}F�(B���)`�I�`[���+E7�!��p�&M��AB������'FjN�*3'	I����p7k���D�-<��W�j�O�P��"����dE����G�7m�#a/��Ӡ�����q(X&�-{������/$���x����:I^�(�g���6�`L����0���Q0�����"��!�Ø̇�3���1��Ƽ�0N����S��^j�-�^i�0-�b���77i7�u�r��T޽I� � �h�& �v-�wQ%o�
8=���w��:
�>����FxEW�|\ba�e��&���
�������i�/��"��2.Yq���Dd*Z��zu?��v���m�u��3��8ER,��B&W�&f��Qm�c@�BD-r|��6�kJ/d�&��ڲ�����jLJ(�$���fW�'j���2���ޜ_&�p��B�џ^��Ƽh��ً�������m�����EL�Sm������ґ�A�?�B+�8g`�g2.<��怍�o�h,b]��=�.?�ܭ��4�!O�\��l�K�ik���_�L	�4t��|�.j���R �4�m;	?��Bm�&�o&��2��Zk��D��[��D5��sE��;'�1��a*��	���⾢ y̚�Hj1�9+�4[(|z&�b9bu���!��SX�P0қ����"=��y럣6'vM�K��Z_�a�6��uDv�͑�v$q�;����p�p~�|'��b�d ԯ&�e��[Y_�jL�@J��^Y�?�ǖ� �T�V���u3�Qey�lQ��E/�Uϵ� ��ZV����#���d���?�E�F�tH`3�W�+E'���EH�o�`�auȊfZ�"�=�'�Y���
�|�;���=�v^Y���<p�`���U_\������*I/H�`we��\�{fb��+�Mw�yt�r$!����[#Y�E�ib�:��a�i������C��O/���~�m��A�S?��b}h<��Lg,c�~BR(���`1���g=+�rv�}4����<1���6n]�烡O����yj�{3���3	?n��"Ku=�g<�#3K��j[u���`��2��ӱ�����'s�ʞ_̤�%�00Fbs$R��S�Xwd	���O-�����������Ŧ� 
�������b*��E��!G|~.�路ޣ�� !�.��R�wV^ɖ��`nj�[��q¥�m��	/C�{�.����̤{=M�:��;y���1m4�R��Juvs,�-���R@�ҹuN��5mɒ�k�bM�֨#�J����!�VB�;|M�
a;�S�W(���,Aǋ#�-��@3ؒA(ԟ(����E�d;�M�#ơ�"m��d���q��G��;��?eX\�ו�.2���tt��܄��Ė��O����y����ea��Whx��tJ �f�GgIZڸH�Ȇ�Y*v�X_�A/7�E�}� YH;D��7h�Ip�>���|�ػ��m�QaW�e���|d�]� h���4�	�dSS	fZ ��H��|�C�T��]���q(F/q>F�E���>�{Q��- gf'M�բ��[ .��`sE/8��#�@z�mU%5�F�?�9���rV����| �J�<�u�'��f���WU��>&y�]�9�b�>�?���< &�v*����a>����0l��FՊ��$����X[ڜ_4�ĉ0U�3�{��c�lJF`�/J�Uh�صM�%���`�]N�Ğq>�_�[���kcM�L
�In�r��"b��Nn��I�����!��T���۪Ui`���K.!�9l�Vi�K��Ջ�H�?&ʅ��
R�TUu�P����å�K���u�}�����Z���\���`�Mpۥs����؃Q�T��'�9��/
�Y�P�.%�@�D��_�1����RC�ǘ<V1S�7��B��c�9�v��K�i��j%�����@7���(�1�3�f����#��V�0�rG�c��O>̯�@D�����dpĩ5��,)�cG�'�^n$�x$���T�ׁ��	^+B{'�3e��e@��!�'hI.�Y�iU��ܩ��֡/�ncŻ��7�I�J�JZ��� �8�2�ҭiƊ��ƙ	ߵe 5<�������'������gN�/A� �{<�lU�i�zA"0�"��a�� �M��� �P)�\�h,���%�c��:{�i�ݠ[�xZ:���&��KL�~>���t�|�O��[״(4T���t4�t;�Em�D���@">����f���K޶\�<�%^����ֺR�(v������Jv��F�K�e�m�Q�z$�r-�ZĖrЫ�O�}�"1�ē����>�n�E� )5g��a*�۽����h������@垢 �;��յ�_����T�A�V�k���o�&m#s�#FT��j��4�"l�SS�+�4���[q|���
�D���y �
b�K����ȬM=%~y�}��TƠ���X���H��2���j����
�a��u��NBcIg��;졝tw��+_��x����}�CrΝ��Z��C�-t����C_�,�6��߫qZha��?����aҴ�@�8֍�HT\����[^��;��)����i�O0,�u��z`s�be��>�C<y�p��B@\X����OEi����6���Q�<�U�E �ZK���\-9��;Z�(ۜ�jj:����Y,�m�9o8ǥ���s\�]���-�� ��mf�č*g�֡����A������A{�S@N���?��m@m�1�L�X�]>Ƚ���3x`Ԩ��F���֑W�.�ɦ��!�hRce#Y%+���5N״�t�r��� ���2��TE�M�r���-d��byn����{$K=����D�w��i�ʩ�<�w�Rb���H�ϨS�^s��v��'Ҥa�������(�U��e��W�^q[U��hf� � ��>{�eS�pp��wJ1],t�ʍ5��m$쫺K�_�;��J��8�"���l�/��{�h��;�B�๚�6eyYKą�fr�9y2��p(0�b���) �7v�Fh�6���'=���_��X���[4l�]2I
�D��,�ldJ��z�q(l��&�K���h��YYإ�KX���VR�/�K��L��.E��h��O�Q�������־|K3�KVg��$��-�MLb^p�#=��4�V��G�q_,+�ٷ�����K��*'Lu�w{�8hx��o�ػ�,��s�"��
�0_��i��-��&<���e*i�o�®�C�x
�э��Y�HL���W(2�l.���a�vE�*tB}�����]������j�`F�A��}���H�ė(�^��QP+��x�sK=�"A�yR�{��2(~i".�����x.e��ΪR�S�ư�(��x?�J��A�wE&t��o*ś�Js�g��Mn��=�t�e	�拗� ����A����o��qm:�H���i�`���s�&gB��~B�b�V�u��p,��$tO�Y����?˖�\�bS���T1l��\�]2���B���i�"��_���0
��0h��3\L,u���g�f��ݹ
n���rqL;���3x��̎h�������� �@����ۉ�G�3�u��AF�B��ۨE�+Ћ����m�8bᰳ<����c]��Z�9��/�;R� e��x	��"��Sm`��D�N���;OG<OY���	���f��F�/��i���ױP���wq���٘癑�8����˳��=���_��-Qp��o-R�N`7�c�ҭHD@�'#�tڧ��\��.;��!�3jS	�{�;�/��f~j�_C�!I��J���̸ڬ���:B���Td-JV�,��~���Q��In�VĹ���ՌӰ��?�.������?����<Y<!_=���c���u���8j�������X���\N�ȍA���������ƹ}�/��O$���SI�^&��V�ߠq�b�I�l�n�~Tz���A��ξ��&Q�E���G8#3p��-�踚�,�շ.�S�n�$ۻ�kl=i����ۡ!�{�����ǁj��8�Fp���;S�z
@���x�_�(���,XE��F�1���%C`Ǒ��~�{%\T˜R�	*�*8gZ˞�~ǈ���b�j}K���]�`�n���v��,��cU���֐N�父ϛ��R�HHb}��YY�R���\3�-7?������/�x*i���}��Mf��߮�"K� ��v`R���f�'�E'K��!���e�j�E�8�G��q<��@�^..�VWF���2E�"b'��Vk=����kS��0<��3�r���+��%cc�B� ��,&B)�6n5�1��|��{�S�<I�,�]��E����G5���0�_�E�xo�D�|�Y�&�X($v�Lhg�7��l�I9>W�JS�HJ��,Մ�i�(�vtME����"|s� �C�i�0�Mr|�1�N�%�����U�՗����:�F������U�-�>�`O��FS@Upb�
��)2?��� 2r�\�tan6�s ��s�@Z,��M���������w���{R�쑿O좽x��s�G�vf�i�-�*�i���t,y4�����1,��"x��N߯�H��0U[u�=Aw�ᦊ�pR�$�{�ׂ?2�Ou�:��
LZ0]��D�U���b��HK�����?��u`-��������%Λ��������7#<-ϙ�93i3�T邞g����cgn�]N$6�R獬 3���zL	a5�{�
��YE�W��\ay�R7>�I)x?N��~/)�eY��鲱�;���!5���1��GUN�kF���]��8��x8���u?���Aֈ�+Mn��X���4q*�P�����ު*x�s��f�!���V��'��G"6�h�Ȃ䀑&'��H~{�Ae|RƂ����$\��M�%�A���`�6�_�Xlz�N�R���Q�ֹ��·4�맛������Џ	C��5�����(��dWʾJv�^oN�}�ģ��P�{Q�n�������a�y��(���7>km�%�h��d�Mh�����~c���h猧F� ���S�P$7H�fO�����+L˯��G���(7f�q�.�dR��Ck�6*U4(v�KR�r�&_�4N��ظH�򊒈B.�A�Uf�?�Ib�XTx#�c���5u=;T��:r��5�U������S��溜."�iS��a%���}B7N���o:0�?�{{��;EY���K�:��q���(�y�(΄G�a �`k �nϰ��5�~'}c�z:�/���s���_���� � ���}���3�v �%L1���^��3��A��ǒ
��Y~��	e��Ej��+1u�4򽚮��5��Wzկ��� ��dmS�k�Yv1}6 7a�����l+-g.<�D�t�5~͹1�D:v����lV_��Ύ����8Rnf[�����p����JEP/X���b���A?���.U@CZR�Ca&�={�l��T�`�YՐ7 p�ž�H�$b%����j�lA䑻p�(A������kp/�R�l¸��T�`�#�9Dc��Ӎo�닚�I��SV-�Ƨ �eP5!� JQ��6�T��{ɘ��"ӭn��J����,w���{F���6�u���:�`�v�=�%�f���.M�D��>=s�*��FYg��'ڈ[�	�_�
����EH�J�ȗ����b��(�/R��
����G9\�V����U�������Be�x旅)L6l��?g�ˡQ�D�\�r' ��F�Ϝ	�<�;��X�Ͼ8`��V{���E���$ٽ�vM�$�'�Wm�h%R!��|�|�3��9VĢ4@�t$��- 1@#k��]а^\P��ү�����:��������S"g�28�����+;c�Ϩ�^�DxcQ!c�σMB��d1E�����\��Jv��KKI���6'9boS'h��=������w�n��a[�9n�
���C
Sjߎ�j���A�b�AW1�io�;Gm̝T����tޛȋ��-�C�Yq�w���GbZ�j�S�9���lآq��1����I�	��-@w5@�B��0g�z@�eϛ"i��)����̩s�2fsWp���
�<@Y���@����Sb~����-���)�i�Lv9*�&Ik�Yd��2�������7nE7m�<T*��+��]�=�_����UN9��ݦ���Usa�qa�B���6��5 ���H'���Y�W�k3̉����j�w��B�X����#n�]B���/I���(W��#���Y��nR�YXQ��[ߤ�Y9G�5#��\�A4a7��I��ȵ��3����P��R7�?fɳf��5�� �PE�������bJ`�r,d�v�Dnj�Z"U}��K�+2|?��Z�<<�R1(Zq��m���Y�.�8:.�]�O*Ѕ� o0����,r�s���t=�"-D_{
7�2�3����k'f窔��bxUl�8�l���	NZ���h7�I�-a3�0�~L$�	�ni;q)��`&7$ �K���z�]ͷ�)���u���g�X�C��W�S�
Dvr��u���c y/�ꑘyOpL�?����E)�'�;g1yaJ'%�<�����I�wI$��e�c��oP:���]�s�ĵ_>�
7�N��`��٫O>e�Qk�'ą�=���b"��R�ou���j)��:����c]�r�vmj�!@�X�R�����x���Xk=?� mz����YR��H����F�T֙�O[`&׉3H�,>�o�-|A��H=�
���f���d�!��ҸԀF��|�M�c_N�v&���ѱ�<��|Nr1� ����w�|�ՊU^R�Ltl=+P�I�#�]50�d�	U@�'���i����֢����;�T�33�iS�щ�Ӆ!�`'��E��6{��J�~Q,�ߡ���P�6����.�HP.U7a���n�(?�`� آ��^��� {4vO��]ò%� ¡��<ŕ��T�2,w��Wj���#z���[j!ȥ�մJDc.T0�*�6��-�l<w��� ��$��{��<O�+��c��Pc+'�]�VPo���\LY�K�+�ǡ�.N�p�I�"b��:�;���:�ɆP���"�g�y��k롚�ֲD�^KW�*�0Ic�Z�jw���I�����ʶӑRG���ƙ�np)�j8���(��8��D��ܡ��qk!V9�F�E�f��J�J�V��]YD<خ�T�����q�ᤠ���E�X&)�h��>�:c���N���{��+�L�VQ�CjSb��U9�� 3ن�_���{M|�"�e$���몚�������S�N_��sh�S�Yj7]���0^�W�?��@�"�����[�=s�2���k�0C��]�Uɇ+*�����5�kA!��b�N�<���c~���/yWTt��wV��h�R6Lف_�����V�Ԑ�P��Ȫ@�;T2[8����i�swp����&
�-�|_��rCF.��h��-���Saf-)��+���Bϔ��ɛ�eS�{��D29FRҟ쵲j��z΂�p�(�b�I#�I�_i(���/C��P���m5��(i�B��.x⤛,�����nzڲq��D�%�L���&���?\#�V�k����*�Ӗ.�"?9d �����Z�^<�6��j�QG�+�]�#�}XN�~�u �tݺrĨ"�L^)��`���!r}��f��p�dY�G��5�������:�[-�xoBh%��mv�:�R-��xʱE����-��.��;��4���}�B��f�(T�gWV�ӽ�Jnyٙ%��O>H�g�z���M��^����M��3h6b�D�~g���(hU���~d���7�4 ���<4��q�����ZYA�*��,[���Alin�cOzC Y�;�fMz��M5�b���G���?X�#��"�D0G%�pV�9�t[:�������vSA뭲�Bs��+G���1Ks��� 6�w�KљO)�u��� ��RE�7������F����B�R�q.�f��������D_�dc2�zM����3�3(��닭h�]�&�I�q9��r���1�B!��R�YB�l�B�α�=s�B�N�U͟�>U�y����|�a�J�}��i���͕Yw;-&k�xk2e/��~��_T�W��ݴlx��b<�{�w�B?ߴ"ʭ���IM���i>h����;QHCZ���BT�e:út��)|��F�]~L��y�)��0�+���C������J�=��]1;e,�#z�D{{&���  #,�0浰���+ s#P�-"���7�h�Ѱ���OW��՞68��6�66@'xrz���������5PV��'� ��+�=~��fGË 
�E������E7S��S�ے�'�Iϖ٫5��?cv:���ۺc�ط�O��g����{eV_�{���Sv,���;���5���=#W��$!�*�o<&���XF��cSV�o:�&5�yK-�?�s"c���\G��&��I>�x%�<���,Bc��x�˳���|�2����������~-�fQ�I9�/�(��\�|��1t��G�eď���β�ZaU8:� �B�[P�i�(%����FyQ����t�A�H�.���ꁥZ�����Y0/i
ɪ�SJ<�M,���!PA�_�Qs�\6��M'T�� /{8DtFK�FE�>m�Ɩ�g/����v������W��ӞY4���ʁ͵zw�yd���bYK-8ioCV��o�|�7a���B�'��R����].{W���p>�Lb<c,ɾp�B�a+�aҬ�~��y�$��ĉ犍����Mc"�o��,��LDf}jZ�O���j���c^m�>�M.�5��HM�G�)����I�r��`��#2��Q�xs�b��}����[��B���(�0Y��C9���c� �A��0����k��j㦧t	H��ꑑ_����Xn]8��1�mя6�����[��\6�����g�a�~�z�@�^�d�R�0�!$.�ǒ�>.q��*Q�:*;-�n7ћz��5��gK��x�z��
�WZ�K��Fa��f����(��ƅ�2@���<]���\톆�z���3��i��t7*Xiaz���Wʉ�l�s��6-�(E7�>d��P\�iӔ-�Fh��m��rY�0�k7vonagu��p�7�č��η��^��/��ߨL��l�������?�eqcT��j[�Ȉ!m��cE�]Y��M���0���2כ�t~dͰ��������D+�=ͼV��G�>>__�y8�mS{�1���Њҩ�������5���r���W$3��4z�ż �a%�i@S__R�&ZeRl�Ӓ�Gj��0̤�E��S�J�R߲�/���A&À����3=~^?�����R�����IT:���n"z�^��b+j��H��k��k�Z$z(g��_��v��P�y�]�e�����!���[�+~�3�.���3\��}�W}E.��O^I�|L�;;��Pl>L��HFc��		�2��>g���p�����\�\��ٝ�Z�9�[�P
��H#_�?�xP�-z6��/bK��9#��kp8'
�g2�7X�4
�s�B�`��U\��s	#ƕ|�^
k��f�R9��iyXQ-YD����K<lG����yT���gB8�+ U��wW����}�f7S�������.��&ㅺ]y�3=�(��
w$a�Zhຫ�pc|�O��Fz�@Z���5��L�Pj�.���a����7P�$�)5E=u�S_�{�V �p��$R��\c���̱*}?����*"�
�f�ć��ᢷ��6߈��0�]C4���!��7��'㘔ŷ�'�� ~/TE�_��'�F����Iz�Q�?��nR���[��G��-�ñ�����!.-�,�[ek�/Q��ki�Vv7��F6jN����?�ZwG�N^ri�����"+����&{����ey��`��)�CwU�:�ơ(��.g(;&`s� ���U��h����3�g�1��}�5-�׽�9��\E�wI���0R=z�.��ժp��~�����>C��JfL?v�j;u 3D
���m{���ȟ�%�}!�K�!���&lD�"�w�����N�ո˿�?°سz�(������q�n���Y!��;$щ�Nt�>���N�_�}0��Qm��F�}6s��j��Ҍ�fȢ�g��Լn����!Ў
E��ti�d�	?�Z�-�b_}�J�Ґ���6�����$$�YR�m��e��P%UXieX;fh�������v
�Q���Q�[����^٣�T\L�Ka\[�>��{���!A� E�߼����y�@5kN�w��0�x�+�@��@E���[9vT���C֙h�ܛ3O�&�sL7N��9�B�#�dWc���wC��dcpUŦ	��i�Wжۺm}��h�Pb���d�����*�o�+�
;�����U��i���{+�z�*1�8�Q�����Y����i<����u���˚8j����k��O�#�����qM�Vt���=��ߜ}�X �S�zEʊZv�B�3bK	+ ��aI!�"�3x�5D7I���z��Fz"�(�3����N���re��N����K�S�lʡo��劗%�Vs�4��6Ud��/6�f��� �Ւr\��E<ⵠN�������F��رB� �H��xVVҐ���礕��ˮ����*#���{����.�[Q�ŽKK��Τ&����R���a9�Ho��Y�9_f��wŢ�u��'\!�#��)���`�TwXw�i�z>���uN�`���m�M�Z�;�NE:�m7��ۑ�4�A�I�ϸo�~���*#�j�$����sV(@G�/��EY��=�[�\`/?�
�YBy����>	�`@�� �	��������O��{U|,d[]u�����6��OA_�Pc��24Z�)b�Q���Ũ-7�-�?ɝ�x)��D�,��O�?�Aj�f6�(N������[��$ͅ3YPգ��-�˜�h��s[7a����ҩ|��-U�Wzw�;x{^(ޔp�%'|S�"%��]�C�B�`^2��׊M� ��_��wE��+�`�^7٘�,5��惿`�)�;ޔ�k��U�6���4��g�5?���dx�*��"ܴ��fjjKC� ��6f�z�qDL�.��.���r��Ͽ���ll?��}j�%�!�ϭ>��͑ۗ5٘�{D�
���V�*{9Q,c�%%#f��}�����fdc����W�jf̱>찳�r�'�0�PŇ�����H����vO4��W���}IT㗱����ߌ���[0����A���^�����+���ú��=�B�2M;��$Ne��m�>\�C��rz��`�SZ�Ɂ*�kI'�fC_�`��/<(�tOB���m7?��X\���Iַ#�ij��:�8�[h��'��)��`E�.MpiJ2��9}l��zo���1{#�����q�SbyI�7�.�& [�^�5�q���H����I9#!f�=64�c2����Se .S�[�u���\݌��c�ơ�n�>�ڧ=b�6��Ҟ�E
.��Z�o���\S��L�"o�� ������R��{i��t��LY��~��]����%�U����#"���w�y8V7�r(����'ٚo��v5�S�gx�=xm\+�Er������
΍��u�}�ٗ���uyfѯ��T�:�
2K&&�����ҏ���y��
�v�^~�渪���^T�$g��ӄuX��"���	�x+ː�����y\�]6��`5�z���,��Y����q��Y+�}����:��rMO��Y���&�s/�y@��}G����x{
�i�!�5W�C������� ����Y^�1.�e3\Wv��g�#�Nu��kgȒ;6㱰a̾�R��8��k
؆�x��̚�3Wv�W_]]b{��y�7��E��N3�I��Tp��n����s�I�"�Xu {�牤�˷Z�7�ܱD��I
lh̘Դ�O�7gDlfld��t���ՕcK#��e�a��у<y�M�vb�۶$i�o���S��a���ȝbݝ���5w2�F��wF�Ud��{q�o���40䨠��C^99(
e�n}����`��_����0�;�@�<����/�	�>��4U�`8q�Aga�
�E�(E�%~��.�З8ĥ��SAY�h З�@�K$�lSjk�G�L	#�UF}��<�s��l�]��׆������c3� E��23��k6�܆�~_ܜ�C�� �ߺh���p�܀�ؘ���i�
P�a�.6֥��H��B������ƫ��x�+*K�����푌�%�~a�$C��8�\T|���E�bC�!����~JB��g�sw�������b�2�ƽx�jEiB#��<!��T$rg��K�_�x���ϲ��L�ϕ� �2͝�?���7�	��*�yB��^1F�#��x�p�e4���\�~�4�y_���~b�'ȺZ<Z�<�K�J�VM�3���O��rl��!L��_�I��C#&����yʏ_kʴ��i�Cߚ�C=Z ZQG����(���N|�A���h��ӡ�0�ʇ����m=�c8HR f|�q(��X	Cg��֕�.���E�!K
�)r���\Զ�P�/��0�(�*)�hk]���1��g�O�d�&��S	�ӊ���7��w�g���� ��?�vAp'�0��EF+5Xە �=�ў�8��Z��,*���a@W��!���wh9���f`��텯i�W2�bh� مW����֖mR��t�%�!\Z�rS�S��I�&k�N���v�ozY���P�Gm �N�I>ˌK�:�����.�ɶ�5YAޥSM�]k��	{I�H_o����=3+�����J[%>�~_B�r�˖��^yCò�ش�Z'?�h� 1��W���DYT������s�Km�MD"�"�N	�D�tV-K��Rǌc �X������ރ���d���Xw�!��<^�X�i���'��\e��S�Бɲiu��P�y�]�!�x�<�O�Q�d�xm��r�=��h����O��{�sSV�m}ؾO.o	tE�LW}��J��FtpKN�C�l�N_���@3��.�0�>Ç���l\DK�F�^����������,.:��Y@�PA�@l�M���7�m�;:�k�w͇��6#���Nzy��q�-�0�E2H�dw�	Ru��t����[��
�Ŗ�$r�w��5u�se��`���b$��ex�B�����0>nX������d��bV<�o����=�86���$rA׊��<�c�����I�Ju���Ú�u��O����@�`����ڧs_0W�4��"썵�1��~���V��r�)쩚Q	]��վ��I�J�U�� hxP���)e����Y�H�PB��ӌ�X���� h��o�1������"D�8�@Z��j���s���%���ˊ�<�o�����ش�K��5b1���-	���5�K����BGd�t��T�4Ҽs{��jg���^�-6�7�ٌ�/W���Hr�L��VԆ	���*t]jM k18PQ��Lk����WSъ���QJ(��>gro1[��X�7�����!�����dE�q��(�[Bnt:s�bT�n,��u���Ћ;�	��X��$���ŕ��^뷂m�WY�v�u%P�ȼ����D�ϼ���=�d>>�-�`����9�V+��xhN����ؤV'��{���V����,Y���A��!�BH�c��B1v�.�����OA�T��Jr��{Q�-T��;�z��wNŝ�3�$�5m"�GB�����X6�,�ԃ4{�U�!B�yt�C�7�I_��΀�#h;7��U3!`��gɄ{n�~M�p���y�{1���T ~ZV@���53�����j)�����\zْ��~�ׯq��������b���imK��|�O=dn7�Ͱ��C��R�z�t�T�JC|���������3��_U}�T[C�x�Cc���Z�#��"��(8v9�3F�ү��$�s;�0��9ty#{��2� ��i�O������w��wwr��,��Lږ+��kM�([-,�}b	��J��8��W���31M)/[ �L{GA�ͯ�j�9Ob� ^5�X�-[}oup4ta>d�e;�kN�M�qi�])�L�Hb� =�̒@��[ �yW�7�������<�Ϡl�@�k8�S
\)V��M5ӂ:�ۍ�[-���Sm�	<�C̫,��.����o0yST��Lݏ�#\I3�"��Ln��ƪ�$�/��O��
Y��e.!щ�ܽ�1��,C����kzK��3	Qߐ� )E��翦l���W��i�ǚ��8�0۝&��[��Og�/{�g��0
�Ё������A~��v�k�F��`hLŖa-��TCT崺v%�x��X�n��_e�W���.vMU�i�@#)Ъ�;*�,���4��kQ}��r9���H�����5��-�k%F+���2�N���\	t�<27�f�V:U��VkH�v��7(j�n�S�v���V�x�Ck�_���/Gq�	j.
����K�
A���8n>��]|K��L�4�����q�1 ���k͜�řE�W� s�KbF��7�`{�~���Q4�u��I�xB*>~a�NM�������	�S @	$P����#ݧD⡉��ʩ0���r$����o���Z7�Ѡ�v�Yv�˷7�>�W%���6K�	�p>�h7ߨ�q�|˙�]���>�z��Yq%���� k�F��e���\�O���k��"cQ�Qi�>Y%Cn(�d�鋺9�
��r����?�'�f�$��s�\q*_���Z��~KLp�Һ�¯�{�����]W�h�I�۴���CsQ��x��KPC��Fy�:��u'z�G!�Z��E�P]�g.>&�K��\H]�xb�"]{��]T�ɝ1b��g�o*�Z�5�RE��k�R�$��a^�����r�{�v��(*iC4�6WJ5�g��4Y2nc�� \73��syQ���ykG2�L�VA?1E����mt��k��U�+�)Dm�BqpSwX�SR������}�onnb|���置��Q�����@�o:�θ��nϏЇ��� ��z\)K+���oA9Ղs��Ȣ����r��4x,���iaoG��kYj�&�\nt����뱧3"&���}|�Z�z�w����z]� @�,��/��x�#o������G`��k��g���n�hTM�,����d�͇L��A���rh�[jץdB�B`�{s��lùdb�qf
��~��yDן��{�dݒol�ڋ��KV��l#^H%]cb?��j���T�0�fx>X0�L0�/wĶ0�Fơ>�	b�K�E��}�|���(�65���^K#y�O,s���Y����#Ӓ�x2Zb��+��
��|��_��:}�[��U(jq�I
IT7������A����m�r��p��O���G ��>'�"؀��[��o����v��E�M��^��:V��L����|�F�􎮂��\�(d꺨	y�焥O��B)�o�˞�ῂ;��Ƚ%�i�:/��^�+@4�U���ٔi&��y֐v����^��EL�	�h�\Ҿ7��=�{z��~��ӄ�?�V*�d�v:����A\˱�eZ�0б9"�B��g�\�v��`�d����:�"�csE� (���ZE���jLp����ߠ����̆�J��>�����7�@���[Ya,&�%-���k�pҎ75��e��e@z G�Kcs��K�Ea��B,	�-l&/�wɉ��w���K�lV�4D�y�ժv��I��G��=Z4�F���2{B�A��J}Z�LN�7�:�Sa#�>t�\1���p�^���ຜCJ��z��%�z�B���^�뎴�z�W؁����m�D��L��H#�rS�/�2s�ü5ϯaN���m�E�����jD�"��k�A+�)M���E�;ǈB�e�v��,�I���AY�"�t���^IHȧ@���O8����ͼ��0pKȓV7>�_l�c��]�Y��W?d�;���TS���>��mSQ�y�|M����i��NU�8�����Oq� u�9���pc�;��_ce�c\!-S,k�N��P�S�T��p�����6J�B�kri;�� Y�g�x"BP��("���P5�n�\oړ|��Jq~����)95�ZaΟ��~��͊�0jt!V����LK���(}_�|��k���&�?�V]/'xl��G_̴ ���Y�B��؃L���^:#�QS�,r��ˢ�\��,�xƔҧs��:�rnj�\�܉O|��Q��6���ǒ3l��2V�>������;_J��i�h�� �)V^-�����h5XФX��B�E���3|�+�%��B�d���;����t$�!��ao ���< n�
n��}Sl�q#�̖rd�5 �|`&z`���#��>[����0vu�D��3)iz/3d�M.����%��᪖�ڣ,�b?�E[��{��H*>�?�� ������R���(������?�Xmbj��F�s0��Mq7�MBk�Eܵ�Uf�?�������`.S��g��s��2b嚨"АT��2d<�E����*�|&�!���0����ˊ�3+���lgn�ȥ����$Z�r-'+5PU��sF�K5���^��DJf���n���aT�� �S�����J
���D�q'�%�9���.��*�8i����F��?��DN����M�-S/���n6Xh�p����̩ŖM�T�,�	�f ���=h��&tH_��f%�z��&Փ1Ѱ��8��G�{�<�X�	4���t!N�B�+���`�~{�m��/��V6u��d�ȝ���W���#�WS�<jB�p�g�化��=�ػ0�׉��}�g*�=lOR��=9\H���=�$��Hk��.�������A��܊�H$Ѥ���@p���(�M�l3כ�,:�[f�Ǩ����G���%�)��<�y��k���g�Ęf���Ȑ_ `��i��`�O�� ���=~�<r轸R�\�ҹ='�
j�Dy�����&P�&�@smM���T�@T���>�ӃM{�ꫧ��|k�t��뭿	�U�g�9������r�FƦ�~]���g�h$���7���pp�{c�꽂�-���a�ei���d2R\��#�>��:K�ㄊ�`	���Qڑ
3�J[��p�"��_h�<Y��S"�C2��$@BP��<�JM3�]N�,�X.ӬP�����,2q	�KND*�Ú�-�� �)�'�؄�N�?��9�l�[��I���3��^�{�2���ae(�.�C����JR��,�FP˩�x\+�Ņ��H�I�c� �[�1�h2�]�.�tev��\�+Lv��P���P�RF�#�;�M&��$�r�*�{j
�|��R��0��Qn�k�TVi��D(��H�i����"���3���P�ц�EL뼖�A?�u���?�k�-
�Me�L
�����:��M�5�lW�]�b����ٛ�tb�{ja����?ǉ�ٝ��*�J�Љ�Xm� �e�ǖ/�5�.q��L#N�j�H��<���I2�CZ[~0�������ݘu��g��μ�^�#��9&�\���;l?���P�p�ժ1�P	�]M���Ա���X+Rt�_:�eX�3�d[��2�F0l�am�WQ�΂L�`6}c��G
ȑM�]�(%o?==(+i #<�I��^���O
�[��	V&j�n6�������� ����dΰ(ѽ}ԯoG��'�H��E!'���о.��9����s�F(�'�'��`""K]�u�����e,86��VR����џ�Ym8%&���Xr�g��]��ť8"6�$Y��Љ�P�\�������E�T�هj���C �$�;�(Q�æ�)����'�l6����f�b���A� cs_�B\��sר41�p{�ҽ��g��XA���jp���K<y��R͖=�L�?��8����ߺJ��і��ƒ�"��.�\���`�=�9-�^���������� %ȋW�c�p�]�!P�k���cZH�x��ǲ�
�%'��3|���ɠϑɃ�Xj�D�)|�Rf�*�`�� �[�~GZz�yB.@�W۲�^�c�>��S<�����9p+��9�+s˜�&��o#|��^�����h�6��m�6EuY�_
���h����б�����M��Gz�Q����X鼑fAY�dx��Q'T�uq�/�g;�y�I\�����z�ՑV��ol��0A�ǆV3ZX�j[7�s���d��/{_Bˍ�#����m$}67���M�S��Q@-mG,�F�{3A�R�̈���]�B<P�r3��m���8bcU �='��L
��R�,�׌F�%�]ZΚ�z�st�N∿��xR��_�/%=��rN�#�BO3	�Lu�q'KEC�1}�c_���z�7���=!�����<�g# ��߻c�)n�c�o������ "2G�[4��Ũ-�ټ�ya�r������%[�)�a�U��廋;z��'Z��2#�x=�iŇb�dom�V�$��Q��wca�3ZWv�R�ٴV�a%8�7�8�ų�͑_~w}�ǯ��j�9����+�� �Üo�8��;R~Ƶ�� �~� ��\Rb����e�Z�:]3Q�rM�r2u�D���2�G[�^�dAլ�*Y��p,����=���@+ߓb2P�P6�pԌ���0K��1�dF1��GDY��15�֕j��i���?+�-�c/��JD�v�֌��+/^�U�Fx'T�;Nz��C&���%�D�'Kp��ih�0�or"���5� @ZU$�WDGGFR�'�E�)'I"<�� ���c��W�
�c�
�Ư�c}-۶�iE�!��g����N���/�z�Ǻ��ޜ�k��bS  ����tg�j�>��Pv�0~�pB8�_�,$���^��G����M����y�v:�����̕�Vc[��7!ݯ6�b�7�o��FJ�g�K����|�޸Q#��9�\9�qz҅��ƶv��tv^��kW���_�F���']�\ٝ�^YBX��BfxB[W]j��]���J�C "��a��/�1�lI�e��t����{��E>P��X�Z��ţN�T�}��Z%krn8Q��>�����I�~����8�Ppa9٦Z;��:��=�t�����S����}�=W�����0�� �Պ����h�e�X���@��3b5j�nV9FU1����i"�md�UF�{���?�^t|#J �������(gR������^��3�+�v箒�fO�M�=���І�n��%n�H7�H������M-Ff����Y����]\�o�_���w+!^(�m��T�s5�ŭ+0`�m� '�.��&B�v!z����'��Dv�|����8/�)b�z���Rڍw����nF2�C(r��y��
'E�~��c���W<�h5mm���K���Y�CX�Z��V�Z�h�x\�������9kxo���#�廑���9����W;��v�n����"�P`��i��6&Di$D�����D�~��O�!��>�)ƪqςE]�h�;9�ßC�/�Ԥ����%�u�w��Z��n�JƷQ�X�7d��_O��i\8H�%�d�*�͔�\���A*v��� ������]��cM~ME���a�9�a�P�j��E2�Y��;��}>�5h��!��2�y���:�Qa���O��ZxPHN��9F��.V�P�-�`8E���q�^ԃ�F���J�D�6U�!���4�ܮ}o�a��=�>2���t�X9�l���U)/k��J� �M*��s��ii�En���5�����ē�vhDa������Jݲ��Jo�./H�G&��,�fԓ �����O�C+��'���6Z\
�z��E�*!ZO�#ai'�ڃ�]{���bmM�V/8�S^���ClaFW0���H�d����~-�-���Bf6�%VfVk:j �1��9%k�x�1+%<(ߥ�>�e�R늜�m�Z=�Ė��~<��눦���B+�z*yXtg��҇o�;�|��T��	H����*���o���\�v�.��qLn���Y0�=1X��Ѡ:֝( ����I�j5�Qdf��>!w[�����l�73�Śi����j�<���g&�ҵL�"��~���gJ�����N���ƿb0�&>�����-��w7��q�s�X��i4��{�#���NB1{���*?,�~��tW(�2T����P <����8
��U��1li��q=7�eě�p6wO����,_zI3��#vڕ��j%�Y*�4j��n����K�T]�8E�ӽC+��O!=Z�H?���d��/L=2�G�VU������ٯ��E�W�h�7q�]��ENܩ�O�M�7�`#iԢ�lCieS�"p�FV�a_���~�P���b��˲��'���u�`�{��1�X�+>���4{[UO�ɡ/���z!�|z/T��d��aYD[3:y�Z�g�!Z
�%s��ŭT����8��g�ux;�L�O�?k�� �c����Ou㉥ث�િR�����~�(��P�3j�$N"��Q���#y�@&�s3��Ȥg P���.!�'oX�\]�laP]�C���z߅c[��lo�X����o_-Uy	;c��'�C�t\�(��ӑ�^�_yR�DO�FZ��!n��/���sMY��I+S%U��ѻHA��h�i4��=���� C:� ��������ۉ
Dۡ�y�֯�������b���ـ{�A2S�	�'3�*F��ܧA`u��dk�{����p�*����&�w�������O�\,�� �@��o�
�0Wv�Ɲ��7*��=`�����	N�:Oytc�'�7�FhY�G
������;%	���Ao����J�1r�� ;�1)VR�c��	��ߤ]��6��8W�����kݝkn��b#z��{!0�z��I)���]�8S�sHM�vi���#d%v%{A>:I@?bF��/Y	���S�D��f�� �;� ��.��^�!:G�F�����S�A�)ˋ��QN�6�<����_��3��-�,~+ƙϳt�� )����I�� PK��k6}iAg;LZ���I��j�xg�	�y�<k��qȲ��o�"e��uDyYOH�{���
9�_�K��Z�@�g�sLݪN���\�#�5��p����\��<'�@?��gSG͇1��h~�ҖC�d�նd�DH��\��e��A�һ�4ӣ�!���ꬦ(L}�B��Wp"�~�[�����̹�yN�cW���{U/���@�-�i^���#ڊ!�='vK��)��� Bb��h�R�4��j-��QA�<F��2:P�i0�9��$-��:,�_nt�fk�.Z����ص�c5���>s �L�k� ����-�����G$M�.��1"C����.q�p#�J��-5V`�:jU�A��6Z��Z� p\�q"��M��
��N�OF�
^���@�Ƨ�����A�����k�>�:$awL9oN�E9��iz�{l�t.kL�"�nc�e��K�9R��^,]�؎���m1�bdk&R�į@�4�we)��ڰ -RU6:���c����Q�@yn\�
_[������(x�������{Ľ@WgA!GECKl�m�}�ǋy׳��ְ�v�����%Ml+��{�*(�������6s[nS��
�jw;��BezﮦIx�fW&�����O�ɯ6�ܐxB�uL��:�@߷�bIK6?���?[�D	3=�`n��J�K�����h(K������L�q	��=g4*�P�Kȵͩ��xv���~Tڅ@>��>�f����m���f[�}O;�V�f��y#K�:`	:��j�uQGL�ۢ�X%dܰ�ef�$+�V���g���o�%7�~xDr�@̀�H�g�Z?F�nq	��4vK���e�8섟�T��^34^fc��~�ڂ�b��eCh�kt���{��Q�i�js�&�Mh҄Ɛ-(�j�E�iU<�^��@q�f�k����ƥ	D�� �3'_�4$��՟��0�5�pįL����XӺQ@��L�M	�W���	Ч�Ҹ����x��d�6���_��B��v�
�;'P����S���C�=��_������+��c�{m�����\N�U|_-�}/�@� ��:^_R���7VX�<�zm��-��1�T�S�vS��FP*�ʓ}µF�'"��
��[V�|���b�hgz��E�!�I6Kbcсy{M�?�{B1o�|�h�����{���̵�,jZ���������P���Y&
\���&�?�g8v��l���F�C~��X�.�R���,A$�0Y/FV��n&4��biĹ�z��Ώ���%���rd���q�j�����L��xe��~j�ky�6�!�}HM����D?N=�[���/���йsK�΁��lNp�p�eP"�a�[`WW<���KI0�;��M���{26���%�W����GB=����~ظ}n�$&���L�L0��)��dٲ��s5�,=u�Y��x#��&�e^	^^�&{�v+�w^�5���p��Ζ���tFR�ֻ8*�%ʸ��@�C�k���&CN��D�d���]�C���\�}���Z���
��C(��RnI�]��С��%�-���=����c%�R*�!P���y��&�f�U���B���]+gV����QΡ�g���;	S����Z>��Kb��M�N�c��* ��1��u7[�vz��FyT���B�G��������1㨎P3��+��)ϸ�T\n%x��� �W�9�OBp��F��(��A���v�어V����R��6�⁷�Xr�C�<I�����*��2C�ک�b�.��h��Y����|�S1���跉�x� ���v�5�Kf6z���C�I�<���ՙ[,J#N��	W"���;���>xZG=��p���%c�s�{k�ķ���N�����u�9���B����x^���������A$�ɀ1(@�9��JT�?`�W(f��n�	�ӷ�ݻ,..!��?�s�K�ev��TD�Gf�}�NVo����>����R[�F/qEJF�Y�8�s{�ӤݐSO��H�+�*~�O�I�.�ʷ���%�X�E��2�E���3���m�z�NQާJ`��B��y5A>� E$�����^��B�n�ɠ���j5��o�?�J=s{:��/��ɃB�$�ͤ��<�B���^�1)�(�я�ʾ�֮���
(�8�$����[c��H_��V��F��N#1$�iR�gi@6ւ�\���O�-�I�Hw�jU�/��ۖ�� ��M*}L�����Q���:t<|6��8���p�x~�V�T8��PgVy�#���਄g�g�upX��)!|F��39�N�<V0gα�I޽"�5M��������j�s����I��2�������'L�����Y��1�!TJ_ه���� آ�����F�^���� ���T-9��XoRi�X�wq{�1�LE���9�����8 T��7�b���w0bQ��o���j�$�o3� s�H��V$�!�E��bI�vְ4�(�N�����@�ν�nX��� 
��f����q�A���.L�4n�� ���c�O<���`�i ;	�G�n��2.�A�K��xd�����];�hE���ӣb(��y�f���-�(�6� ��D�
M�=��H�,�ڌ���~BM���x/8�U.��B�.���`޲���`��8�2�,���1�5���1��5�ŮBX����p~`� (�w^ǀ�V�.H՚�[��~�-Z>*�S��sA'n��g��R]��崙���O*k�\xw������i���&�.�{ů=6�RCx����9�|��y�L�F�:�x��ؕ�Ϋ�u�u�ώ��|Lh�|�d��T�}�P��I��u)	�C�^��C�N ��2��`߇�}���	�Q��wޯH�P�!4G9���)j:��n�t���g9($�/1i�gW+���8�i,�:'��H�2pnhQTo�5`�g&}����-Ȍ8t��8:�l��(�8��!dgG-�$~�:y�&R�^ˇѷ�X~��eY���@A���5�k��Q��vl#:��ZP���C��l�4X�1"�����{Y�#R��}���1�gͱ��r�ئXh��=1jɷM���塞�#X��e�;EJV����S����9����aK��xf�4,i�&�$ ���"���ּw'n%�S&�ж�V��{ΫEӎ�]�*xtU�Q����`[��?=a�{*�Aeϰ��Yh����R-��g|f��x���V��r�u�u5��7؟v0�s�G��v3���`&�r��L��CC ��)�@�F\�x��ݏ�`gp.f3A��r��Պ�W��]�����hb��`"ae�Yx�Z
������$y��?��\���K�Є}��l58`��Z�/��E>u߉-2?4��; Yc�+�����p���5%&�U��%�sI='�(�.�Y6�z����fwI���,�wÆR��Aݷ�Фv�0�֙�󱓂�Y�nK	%m�iyl��r��� h��.tbb(���Tb5�T��D�X�@%����)h�
��Z�@�g�&|9N���u�[��9��K��`�4��v#@U��V�m��ǩmJ�¯r���=2̞h�{�d�A��5�:*��9={z%�p+�~�*6��L�^�{�OU@�q' ]���9���3��C5�-H���w�Z�!�g '��pF�"d$E���A��_Ny�U)�^��'������Vjp�]Z"�]��+q,9�#�n�j=�@*<	i#��@x�ix.L��>ˢ���:���m<9"���oeG��,H��?�H�Ww���5�dWi�	.�6�����̕�+�PhĎY�ea�/�R�P	���y7n��b��@�����6*j�K����PF�<LK���2�FgG}'���)ud��1�~����O��Hd�/���˽�sZ�T�M�H̨��|�t�%�.��CQ�ϋǶ=)�%�V4S��M����C��؎b�V_�L�+��>�k�H�ȀTb�?C�2pA��a!��q���*��A���A�{S��ҹ�N��h�!����-X�-c<���R���s��i�vl-��c� �)~����y�����lj
�`�� j�З�����/�A���y���r!�F��V��.�jLP�>���gh�vW]RJs����Y�^h���Y$�}��9�g�}�CZF�Tݛ��������`G�ќ���VO3��O��W3-=����6�`d6�"�u��������Ba��&�kb��r����i���ʈ�a��]�Mzz!�	�%-v�Sw~oS��lɱЍ�4G�1�\c$�;[Uް3Q�	"�e��]]���'1њ�d������ު�?&��W���Zny�#
����tR��������ϛ���j1M�U2T����
1$�xlꖡ괙!�l� ֓���*y�xY�֜.�q��ۘQv2����������6�L1-qe��8�?����ڻOE�T	�]�ޣ����!c7>�q�5k��"\�g�B��@�ee��������~��\lh`�bڏ���|=ҡ�z�i�a�)}�0#�fY��X�hJ #�q��~�z��S��o2(Ԯ�$� �nb���Z�&s�� �ϻ�	F�e���$p�
��G!0�����+������D�����@��k���=������ܒ3������JX?!��ԁ?d�1g�'�q�۽s��f�O�۰��;ÏN�1�1��5�\x\e�&8b]�����`됖��m����,Yp�@��N}���V�lVk��9���Ҫ����Ry�&"g���R���ٗ�K��v{ź�O��U����j����m�����6K_\%o�G��!&���p9D�L��*�b�� �D� �#GE@`�ɴ�����đ����կ:���t	U|j}>/�f}c�ͩ�tI���k)?�c����ȳ�m�3�nk�����X���uN�C�n����cw������������/���"i:�>��99���zKٍ{ׄ����|W�¼�C�� �ڂ����MG�H�g��8I�����T�v�1'ҩ����Z;�Юn[x`�w3�Џ)�KH�<P
�50�媠�X/	�~d|�����[%��T���Zh���a��p>�y͋Ԧ�� De:��U:���������ZQ�-��·����₹E�X~�%�?XH�9�^&��>�@Rb�٭|<fb8�Ga[����i�����}@'jj-�H��U�3G�(	�7{F����)�<�+��4=�g�E#ƒ�iT~:=�c���T��p�Y�.���^Ek�a��]�b�T�d����zJ.ڜ֍Ɖ����mws�>�cY�Z���i�t 6�b��L�'�A��ߦ5���uRl	MOJWadQ]e�0�P�s��퉒�����KAw�mCG�y��$��=�;?O��;�T����Z1lة��������2�8 ET[�u��K[re�?"y��%�,�&�����9O�Δ�הּ��ٯ�/b��s3u��So�����!�5�`��34�{nt���J�K[s��gTHR�4cGH]�L=�5���i������0g���W���U�C��%�fC\V��p���:.%P��pA���n��D��tO�hRa$��@�Z%Q�j�%�9<g��DB2��Q�~�W]���=�p�����C7V�~|�̼��G��ѳ��6�i��Ϣ�7��RG�?��	���E��iV�a�g�����nq�E�e�̽P�;(���x4�6��D�۲l�Z���
�Q~�+���o�~�4�3�.�LBI9�
�B�.��3����zo*�{����̨�H�?96��Y�����o�)ROu|��#a�3Ȗލ#b'�3r��%��/�C�@s��o�i��'�Q�t`{%X��u|K�!��9X=j�$���mu��(�iGt�L��on�Ɗ]5�7{^g�!�	�% �Į���v=��xp�<�J�Ao
����M�yb7�[�Fl4w���35�5+}��
4Hj��Y9��0�\��C��ί�;��R�t^���Q�{���%�d��M82��[C��r��yO|�]�'ov�`	��o�`�R����S�w�=U�/�`�Z��Wx�0�uVO��HZ������}%�c�.~�߫�+JXt�>jU>��W������\���WNA�vw��,�K+�$��ܛ��>_�1mV�3l+�:�yk�v���O�ME���Z�8_�,��d=��_|2i!#~QVx���I甇����P�bF~T�lRf`�_�}#v�C��>����WMTX�4ď�#� ��^���&x��v�ʉ�k�2�=ޤ�h����HnY��'K�q(��K�"�I�؝��ԗ�N��M�*��������)�l�Ym�!�!�E�~u�����fa��7�R����G_2����W�F`<W`��!r��`y:p�'ӫ8�	����Մ�зĠ�JE��	���RL����*,���8A���g������+O!`?r�/g���3���~�adY*�$�%��:�I4����|������q��m���;�2���]�=�Y8��2Mp�:��D$Q_�"%�㾫�uD4�	���-j��Ԗ(gӢ8�f�i��ny��c�z�;!Ʃ�������i���u6C
��Q�0� a�ދ���ӍM�ܐJ�d�~��*x��}���o��w��i>X�q�k��O�7�t ����{`�A��X��<���|e�v��%����Z�%��{M��i�k3��>\��s�Oѐ 9�i3��F^�m�?�����A���Lg�b��W�r=;�l�8 Nf�ò``��S�)���Aٛ�-`��a��݇�v��RT����\4�H���K��0bJr�CH_���J害 -X*'�f�0�	��/GYg��f�����B��I�X���L<�*�6��·/��b�7	z�Ϻ��W�x&���:���)���;X��
�4O�p<H$ԙ߄)��55:����W��%t�����R��ɓ �ڻJ���^�0�1���g?x�k6?<�� �
>�S�y�A�z<�f�DcT;��%��\W����0��_�;Kc�%�{��jPp�2�.�z����W�D�m��)��`ꨮ�Ӛ����h}�;y�)��w���@?!F�!��8�(?=�\\V�7Ȥh'c�	�yb&Rϳ�H��t*۬�
4"���hV�'D��[�Y�dqy oJ����,T��T���X�D�m&{�+���ѽ��&��$͋�T�g�[�3W+�TMm�K'�wu��QXw�h��'g���Оs��L&s��XU4K&Wê��.������u[���]��f�#zn�F�A�+�_���:��Zma7��b�ͮ�7�o4��9��ˎO"`�y��.s�_�;Vp��J��-$��cNmh��u����	�c���¦tg�%=����g��F�,N^0���3[d�nR�5�F�*
$�<u�6��gI.0����eH�rs��4�P��S�1�ܮ@c4V2f""Ŭ,�)��s+W�L�)�$յ���>�硰Q,�c'~`�Cx���5�;!K�\2QL4H"���Y�>�Ҵ��JR%���xKjC�YI�[$wu�"2^3g�9�W(�������ㄍ	+	4�x�� �2ل�ą��O_�G�<��,E�d���%p
���K����Ц"�Z��
��閘iYב�����TPV�l9IS������$_}=_���]�`���G�ȹ���ׄ��$��Y����^�X�L���?��O�:����B������j�����7�C��%@w�]7$��7��`���S�CK��~�����Ps�Wr��*��uo�R%�d��� ����[�?yE�����Y7]�5ݭd}��=�	Y��O^>b�J�k[�:��Z���~���r��*>�';g�c�W������"��S���������.a��~i�`1��4�EFc`,�bj���bft}��Ѯ9 O�.&G�b�<�O3�����(�q���$��m���Y���F��Y1�QZ��X�;{KI1ِ��6/ܥ����
�4��D��b��S�~Krcw_X�:Ǟ	{�>���Zi#��sK��P��:iJ�F�M����+�Y�%H �{�V�	�A��~�}���K�5v��+N�--�%mv@����󈰾.jkh����6b��X��O7��#��#_�JS�+� -Y5R�׍�������4N�m�-���c�.�k��\a�!�7�=�Ɣ3Z��w'D�@����d����G��i�v�a��8�8Wq}��.�r/�9Q�'��̢�Z��P���⪩¦����v'�1E�EW��
��_{�S��Mv֢�\��(��5��(4L�g@��p�( #���C���e��E2��e�ߎ��Z]C��0^w�%�	�y8���k�}�y҈�����63��Ԕy�i���96�.ҙ?{|�wb$�)o�g�|���9>��-�R'�ޠ���J�R��DN%�Ds{��!�Q�a�_���8]���������c�P���{�o܁^��(
o�Ml��.�Y1٥h������SO>������M�`1i�>�VX�jDN��W�a��R������rm�`�`���{��>�Պ
"�F��r�Dx��/>k.	lI�h�7ؾ�}����".t�,ɣl.`���GlĜ���>/����0j���xna����T@Y��2ޱ���.�iP�;
N���Ah{��{�v�H�U���Ϋ�IW�5��uw���ښ������I颮�7*����h�Y�ei$����l��}�rn5%�Fa�#��O�_u�k����?QSa�س*b`����-W�L�f�u0��`f�ܓ���V�I�����¿�OcgY,׊�$N���,����(��t�g���h�m�ƞ�PA�Q��Z}�z�"�BJp�s0�U52����^%h���P`ŁQQ�����80n�o�0�p"m}�ճ�B���#@H0>�iw��y�0�=�K��Ei��`J�LkƏ�&���`�*�턫��&/SP^�m�{M���MK�!a +��/���+L�F��]kѳ1eXO7�%~��d]*s�PB��/�U!!����IE��0������My0ؘ���ʩ����$���;�v�v��Y�����3��v���U�=�<Y��%Nx/��6~�ԕ.�Jb@�8��A�P/~1��>��4�z �XJ4���ʙ�j9<�8�z�+�R{|6�04�ܦ�Δ1��}�o�Q�ˢ�L����N��U��i�c��H^z/V߇��`G֧�z4J�2�-3�������E7OG.�m�O�wWy�<^�2l���y{��1\�j���T�kvp����K��h�@�Z����o[��*z�����3C���-? ��)F4!Ip�YdяÇ��('��zx<�ˈ;�P�g�()B=�V{$u}�.�]k'A�f�+7�P���#}|U���Ɇ��#fTM��"�i�����Bkr]�\Ϲ"�Q����/�"�y�K��WX<P�t��+U(��9�MO�)ժ�ͩTkGE@�7��Ax�5�t���k|~��&i:[�������}z_��%��|Ѐ޽��(�L�a�V�(�CG�{��nO�b�ⳗ9.�:ݝx+Hyer(�6�.��f\�R4����) Cڤum�c�r�����<J�{@���.�aL�I���������'����-�ww�sQ�C6��W�6�oT'��_.��t~H����z�+8P��.6�ռt�l��H�B���)7�%A�9v)� Yun�;�7>seCJ0 o�0���Z b�V-�h�\���Y��x ,6L�k9]�{�'������RjO*5��W����K�d��֚�Ae����C�����f������T)��.
����;�[=�lA���Ă���5����͚��5�7ٕo�6���3~�w��gci�=�N���������ŏ%ҚrH�:�HTʅj~44�rM2q ;�}�'ѥ}:t%��Aš.�5��!)焑�5ur`+��"U
ۏ�wQܭE�\�Y`�����,���Мe��X�|5?2���?�����-�5�;��A��^�߱���+|>c��|R%���Y�Kc����X��xӚ��\0���z&�����7|��?(�x�����ZRr��l�؊>����z��hSn�>�@[sb�  Ŋ�/(``9i�4	?���Epe':bw�"�X�q��qW;�-C�)74<&�Z躎kmԗg���P�X�v��pչ�Bm����ݷ��]h�6�{� [��%��f�rQ�r֭�J1X����n�1-��8��r�Y�U�iI�2�5M+-,��!�(�j�͂'��n��\�E����SV�y�ʗ�j�H֠�e-w_BY��og�[�Q;�9}�D����{.˳����n��ϩ{�<8 }��ѡ˵ݪ��:k&c�j��|s0�� `l{f>�f�Η����@d��F��l��HXS�#c�آ��H0"���FG�
��4Ó�ڮ�o�άC���ƪ_��v��n���^ �*{-�asZ�u�=I�b˗8�����m���EΙӘG�)!�U��WX�Y��"�,�eas��o���N�!�]]OD��n2D43�2�$��Q�B����a�DvQ��h�����*ٷHe8yB�	�W�E��6S�y���ϑm�nj�I��2k� ��Rr�(�0��\`�^(���^�#������'(I�k|����q�f���?p�g� �2���9�bv��ކ��a���T��EO�'J}L��+����",���?��U�oq"9���ye���CG`����z9��w ��%:8��Z�i���F��-�v}�v�GD�l��e�(����F�_1T}B��N�ч����p�8J�`�~E�c�mנ��}d��.�o*�=��B�n0�'�b�Qu�7�Ȃ#؈lP��B�SC�q��X~�$�e��$� .?{����Yׂɞ9ҋ��<�vd���"$Yɪ���Ω�,BS)��:�?�T��w�J�ЙU�j������#�2v���@R�@]�|O��O�R��.B��E?@9��3�`�a	��oU9w���׋��T̚�cd��?H%
�j�k���+Wq�[���D�ڎ��{�4����_0�>�o�ˑ���W}��0N�q����t}|����[J���"o�h�Pԙ��c�#��[4"�K���Y���ü�ʨG�6��&�wl�k��PE�8�0Dt�3�kx���AМ�6�-�X�_o�8,���FP﫦�;^�Fp�i�˟y���c�Jx�w������[��9��m�@p3�������2��+��#fU�#j���jfh���}OpMV� p������2���g��M����_�QDk	�g�6U��{N�]ܨH� ���zli�j����uE,�i��9�lt!lŢ��?s��3��䯑 +81UW7f�[3���s�o�S�O1�\�^�o��%<}�\�����!Ԉ�|uw��>,����d�Ey�ήR{��&�-�<�l�&a"���-7��߹��0jKQc�0�M	f�+^�]����'�X���3��m������A �JT.A*|kW�#E���6KV?�����O�c�8�9���Yh�_�6�m%���d��� ���Z���qS�Ñ9��ub��
\gMF��c����@|�����{�z�M��䝬"���4Ӆ8�K'�M���L�5��}|��c#t�6�S	�R�b�\�裿j��s��d<,P|�O�]����
��+W>n���Q�P�5 ���V~��qh�4�_w I��)��i�Au��� ��=�B-�}VFO?J*4NN8R�\��&�w0aS��z�Fr�툹�T����:t�C4*�D�~`��	�A2�琈	��m.�V�����TB���y��'�׺$�r�?v{�kv�쥘�b
�=���|�Y~rXb(!�?B�I�k�r�"�M]�w�����5M��4�?�k���`����,̐i�UϨ�#*}�Y��Gٗ�qG�qj3���Ll�!��2u��S�^Y���z�J��B�)�;�p�s��z^(	���5M,V�	�\�`p3�	/l�F�/���ȧGġ+D��Ƣ�u=c�5v(����"aj/e	v�c�	�|���ľ�({�ˈZӬ�e�m�F,5{��CΦ^Ы\s|�$�����F���]����#�(�$��Ƣ��"'�p��v�������6~���^�D`��c|�줎�As8��j�P������Wˮ��XC�	�`QX3
0���q�&PUJ,�+���ֻ��k�VN��H�?|lKU s�{��Rm	s"!�h�o��Cl̾7�-�B�TN������
��k���>��v�Pa���N��-�Y ����+s�Xw�
D0*&~_!�\��K���>������˓��W�\����*�DB�GqV1�d�b}���
�;���F|��_p_6,�i����b���S����[���oDO����p稦܅=�k�[�*�����F�7n���v*]�W��g2C����Ê���λ����n�9>WC��8�}Wrf�,X����{���cem�c�N)�L��'S�^��3�q��g|H۵T<�4�1VOh#x|Xw��i��p��g���i1�����I�q�L���5C��'�9�;���[���.Sː�L]�	lx���hu�g��NQ��B<�c�(J4�ѹ�{��g���~�o,z!3�S�?�R���
.T�0��?�)b=R� p�_�PQo�42Ls�_�HK����Օ�X<B(�\(�	�kfj���~~C����b�/�O�Ƕ��x��H��|%\�ڮ�U��6-���D9�/]�Kخ��Z�֞�z�v�C��&*bF0S�8��2��fyâ���|�b�ECp�����G���,^W�������@�=+#���Ͼ4��)�r^�g5b�L�1m^v���َ>���w���/	ѹ�?2�	��ȇj�m�>��1���5��)�^�e���1*� �J|8��ٞ&�.b���>P����� �~�V���3�{T*�I
��;�s9 F����c�������v�4��Y)S���f�\���ȹ�"e%���b�������M�H��z
 ��vX������yt������n�-Ji)'�=D N@��R�&���,N8����Sc@x����W:���P"�mm��6�r$TLEl�/��p����B<�l����I�X?)s��ꐼ�҉�o!/-ހ���"�vEFs�3B~*Je�F�^|q�֬�'��z��OG�g��X�:#�ȷXg�Bs �n@Ɉ�����@�t��QiN�c�[3��2�22.})���o���X�q�2X�S���3gx��3cL��PT�� B�܁tԫ^��K���]��Ϧ��F���6�8*�N3�T-�Ɣy!�;U�&���5(T�%\dwm�IfY��.�o�IM1��o{Ĝ�fZ&2��݋�_�<Q9�38h�ƒì�Cy���I"���^�ʹ�E~��/8IO@�o�;)��G�{'� 7M;��`��N8C�U���s
�iC��zk���X]|C+����:��s�z�f*��h��͍4��+_�f: �	�&6h�a|Jj�J��ȳ;XZ���=ܹ]�W:��|V�pQ�Q��^�HV�>�TV6�������t�lXi���J�����E�/)8���N��p�U�.���TN��?l��1�tp1'���w�����M�<k(�R�5ߡP��-Dz@,82��{�+6��w�'r�C��c����� �n��[nVPe��-�@J����ݖ���F,�m5��U^>7��Ah��Ah�W�������U�W��^D�1��?�>쑶�`_ȕ`����60��\ǥ��J[�-rT��ܲ}�{&�Nh;pN��W�Lm��l�&}�I��Th�h�\���B�6oͬ�E3�GD�ـ&�`�9���o�.�j��3^��������6�Q�$�����$�蠄�{��V�u����ظQ��A$�=� �r�Ѭn ��ڽ�=�8�~����
�
�XQ��,5y��k�5&�3Q*3�4!X3]��0�%��c�1���)�j<�z{`���
'�9}Q_E���q���
؍$��`T�z�B� i _���_���9���gj7t��b/ε"������8�m���=�����MŴ�|�A����B|�P !����k���Q���s�)��l�H��;|��;P�dӢ>���c��֠����|�U�x9<�Mm�(���(��s%�͌�w,xi|(�b .��y��]�v�h�SA�����:gl'��1��o�`G��e�@�/l	V��I+�j�̈́���;����{^qɤ��Y	!bD��e��{���jiCP�o���CP(�����+��d���y�RἷO�{�X�ږ������ߍ��ƴJ�����@����=�NK�~d�óS̑���cd��pX�[���Ƀ�8Z�������{!fu'�6�k��W�ưj(�"Re��W���Q�9T�%���
���or��*�-��y�3��(�[*d�ŉa��12y��nB�R�8"��� o>��)f���Hb�J]�/�[ZX	��j��5H8�ԋK7���)ŀ����ͯč(�:��E4��3����cɼ,��}d��u�l�^ɉ�0���5I�i.3��<����*_+Å;��Q���*�薚��������DuL�"A�{Z��6� ��� ?԰L[ӗ�Lۏ�eC�bR���%��Yȁ���a6�39�Ƴ�$o�7T�U_j�U3�<�V�rl��Gil��DLv �%�2�R��o�%���$4�<�T�*�_0�[8�z�o��&J��
�R���~g���`�+����{��Z�6M��Yq�+F�mʬ+G�j��=�&fc2'/6\�k�Ź'^��u���Ep���Փ�mm�F9���m�a[��*Fo�}J_�ݺ �^�x���g��`J�+��o�[@�m��ð�o�*دmÉ|�����@�c�r�z|��ֱ��@�(Q�3��h��yj�[`��H[��&a�~#�䞮i���f=�{�F,���r��X��ś���6��LO�U�ꪡ�9t#5�=�lO'�}3*����#֟$��|`$W\4��y�Dw�aK���[E�DX*���n߽C�I`΅�_�V���F:w�e_ͱr/�ň-�+9�3����%��	�$K�҄4�L%���w�����i�R��/'qU����/�UR�ĉ�mU���5�zTufcI����&ngd�hI�ekΩ���&'�y��I��~辙#�	O��ݰ�e0x��R'���5�.�ds�k"~R:��Z8�Z��~AQ'���er�>�$�r�u��W�����r���MA�o�X)x\�=�>����L�Y��X���vF���PTH���SeXv��W��2y�t�М������o��S��h�K��/W�ԕ���w����)�����0��d��c�$9�Z�8��5��������8~�#�]�wN��{<!������[�E�\t�~����"!�1����^�HK	��6dg��X���|�� �6d��S�p/f	�7�E�`G<��k�����)Nx�D��>��iVW��ٖ߀��)���zZp'/���^��I��z0�=,�L��,W���.*xE���]��f�v�N"�����T�g�hz@�i��&�fv��c}K�T���`���'|�+;�%M^]�+�ro��2�f@��6��Bz�]0j��A>�+�B���������������8�3�NeE�I�V� ��q�Ѿ+�]B�p�Џ��I͗N7�X�fw�?����Ū�I	J$o�Q+MB�кTez���6���;�@s��O� �	kW�j�Gt��ʺ/���R�l ���oS�4.��ji�XG��M�x�LV�)D6U�W�|�q׹8ᖂ}:�X�_�U�aʐ��]�����X7�07�N)#�p̿{��;]�(�z��]C��1V种ۑ�x���{^��K�R����DhK��I,&@����S6-��L\���f�W�|�*>1��w����V8�r")�V&q���_@m�j?���2v������V�^�|	ug_�H�'�}��#3��GS����}p\�?�M��=RnE
1�$$\��<]wFB�]d�����SL�N�����a�7�g�,�I���RD^4^�F'���r%⹜JW-���$��㲨��Wko^�ڄ���\�2�i�w���'6!�Ђ��֭��H����f�	A�%s��ug
����}l�:�`m�X�]���
���7}AS�e�c���>�/<Z���sn��,i5c�M&8�Z�G�U���$�܎	�xp�@�M�/��؏I<x��K�s YRF����qx�3ry�AFM�tZ���ѓ�oE�n�-A�W����=o}����ur$�@��n6:���z� C���@�����c�J�vd�psO�LZ8ˋ+�!u����g�� �w
�W�]vf%�Sr���?o,�
�bs��j�Ov���vJ�>�����GhH���y�o�a�.0���I�N��Qs)��SG	�:���z��渰����!װ=3�ǭo�N09��nE��r'��4���*�}��
a{�x�v���|	yC�)2�U���z�>*آz���J�B�Ͱ1FH�PY�����vNv �.��Cӳ�4�F�K��f�8ӄ��l���M�Y�Q٫�Ƨ�A&���'�Z���:p$Xc�n��m�����;W&v.)��y��{�=Ƌփ���a�+̷�rqݮ�.s��w�&��(&f 䇥6(�8�f�PC#%��2Z�w��Y(����n<�W�����\{�[\]4�D�1�n��7�н�G�B�c��w�)�.4��O�S��j�"&���r��E=H��Cv����#%A�B��,3�p�����$&�*��ߌ���t75��)[����bI�y�HІ>��� ��	��քO��e
�aX	�E2�rNn�>,�W�Q���z��,b	vC\C��s����u�T6���c^g�R�dT��������r�����	#ވW�x���Y������d9.,+��M������z&d�tT_����x�Z�2�zq�c�.g��%x:_��DU��t�S8E�U0$oW�I�rGɪ�)�@w���}>�p���wK��[�D- }�y�f���<��w;�+�k�� T�AЄ�d$�d��mn�)/�/�Z�%<nVX����H��`
M�3��gʶƎ=f>*h�&��lg�7c��B�\>~i3�d��?�))c]�����5���TP0^s���ɠ��~kI�*o+]�B��-�������6Ur�g$7���J��_��vy�\f�w"M���!�o�D���}Gїݰ�E��uS�������\����D���"B�=a�w}7����~0�Kd_y�?y�c������"46�Á�_h#9R�"H���t�D�m�м�� ���@Y�Ǩ/i���aS��2�EQ��.�������5D~;/���A�!��=�Gv��,��e�\Gf#�q�[ȻG�0����l��������|�W���{ְ��N��_���$FL[,��{ޒՖ��P��ӥ.oD{ʅ����tB\�:ƛ]���؆�m���H$��v`톮�%Ez[�|UcHI`��pn�������4!�6<舞��G�[�1��i�c�拍����xG��yC`e�^�.����a@z�C\�~�=bނJ�{�\}@��E�����͎���^$Yݦfr��>�m�O�d��w��q�!�h�M�Ü�m�ˠ����T��Oo>�,����O���K~<����uE�;Cs,�n(}�R��D�����$Oij��f9 i���UI��B��˱�9����+�PF�ܽ;�(���vD�El�\�qCJ��C�����c��Y�8��ކ�Y����W���f�	���T���cTds\��ru
�/�˕�]����&��/Ay�~d6�",!���^�����?I�C&���xMJ/�K-(KK�I��^/.�8H#��l�-�g&\ڔ�6��X#���j�r����W�I:_��Uv6>�s���R@���SV��<H�胆���J�����{�7���*�(�9�?T$:(_:Δ�ϕDX����A���\�jӮ�����]h��,WX[�4T�7E2tw�h��{
 ��~���  `�J�4�3�!���F����4}�i�{�k��\�������}OwKM������Qm���,�v�����MI�j.Q%|�yf��w�,M�o���D������ *�"�UVs��#�X�ީ�� �M+_�;��~\:�5��0�d�
g�G��{
��Y5q0�Be ���MrF�XB�@��|3��K̆V��z�����F,Ng�ӱW0M�،H�ߊ\}&���<Rt��3����lJ�A����5�����u�]�XrF3���^V�F0�� ��2�ؤ�� <A��23D|�R����Mxi����^{�l�5�����b��
�[G�~�R�䬔0T��A��[R�Կ�U�p�1��S`灠>V��6K>�绪�N��M��(5u�1C�a�{���2*v�3տ
dp��bvN����K��}?U�k�xǚ��ԛw[�b�p
Ѓ�ڑZ~>�2k��NL�Iے�s�s�u�z�]%�}�`?�b*���k+�qVyZ�.��@���z��IY�JuR�����OP�l�@(��@{��Z��cQ�f˨cJ��f�֊�$���	ϵ]��]�Ϧ5�3��O��o���fS+��v�?DG���іRЄQM�C;�p�h�(
�_m[p\��:ƒ+'&��T9��	� F�Jo8�B��oG�d�'���Z�S,ZEf'sc��&}}\��&5����=ڈ�yf��|���%,dmV�[���ys"�w������i.u�Q˿���K!���.�qV�ԕ�0���&���xz]�e|��[)�6�1_�E	#�KW(s��{��6�.���6�W�K����}^���*w8�Q=��Ɉ��R���BO?�k��3Q��8����黣�v�GX�1� �G�?��H�_9�y���Si�'�҂_��u��eg�ՠ �z���X1C^��7�������{a��k����؃���F���x;(�zw�k���LK_+(1�G	����"��E��oB���/�< ��.3Gy��SvGƼ�ʰ~�Ϭ����f��Ʒ��-� ��$	`Ew���S[��b��~y�
�"�T_��-Ǧ֧�ٟq���b�q12�_��1��6�uA((�cN�+\�9	���=�-�BS�Ɍ�M8F�O��❺9Q�i��Ȇ(B��[������n�V�����,��K�����P�1O��(1�N�Z�`6��h�<pUD��k�_�R|}�8T�|$�v� ��if~��h5�.��c,�OG�E-o�`j�e(���̦E�	�:zw��i��;��/�g8U~����P���c\%������D>�~�hB������{!�|@cDF�PU8%[=�mJ��8��N{[W1��R.�[5�	�����^��|���f���\R���DW�Y��{���4��M��k\��C��8�	�A�`��nP:����H\�;B����F�̍��?2�{�Ņ:��h���VY��a<�,��p{w'n]��[-�l���W����f)7n�X�>��ǄfY���7�֘���Zs>��?uT����s�j�2�X�țB]t��Pf[e��=�-&＾�iZb�u��f\4��O
`= �3��]�k�ޜO�4�|����G!��z7K��G�6b�x*����'�V�u'3��^�@�7�杤��E��<*��rDA�"�s���(�N���D�����va���9(��vsO�a�i�?De�����n�p6���j!+R-��� Wy[ƲH׋�����|Ȃ��t&�K-�oD��],G���A�
8Z��CC�a�D`�:��R?�@H̨l�(���GO��XW/�d }�l�D�K؍�=r~�Z+��Ib��2�Œqy��+�)��4�u�"���5�"Ivk/P��n�OlE[\�&�PƆ�������h�~4����U7����w%G�ݳ/�b�c������S
��f�2)豉5��,���EW�� �\O6I���g� �[
?��{3�Y�(��2��@�LԊ^?OV�X�z݅.�7�᫧�4�.� �������å5�dC�،@6�B_n�d�A�s�9Ǥ�PK��ՙ�k���u"Iwv�&�Ѝ*�K��	`�g*���bf��c��v��1�h�&pb�:4;|����)��"d�l���%��ַ���M�G[�X����e�d���(r��I-�}��Y��q� �\f��?��/FR6��b�(N%�'�?�(�������!�T���]d��D��5؋T]�( �"Olݯ
r����~��1�Vh3� ���u%(��
�Oc���n�'�BS�(y"8���J?��O��'U��� ����LМ=,�gL�#�@�O_�˨䞰��Ȓ���!C���r�±c�B(����:�Th�U��C�"��?�|�˼:�<{�?�@��M	�t�ji+�%-�W��x]���� �%�;Z������(�:�j�@��,K�%`��.�!s�!�Q(B*���4�|��#v]Xy�b��@��e��u��8�w�u��8�˅OW԰�ݗ0gҢ��q�|���/����VG�a&E��*Zm�D�s�[]��g�V����Bac��T��m��YF����*�cqCԩ-n�dV$�����,��W5�	9}��Q��D����H�N�,L�H��k�.�sV���u9U��G����.~Q�-�c�v��5M�+�i�:3�H�nT�c��z�|[��m-��%~�r���$"��OTþ;j��J}h�aД@X��������)|t�!�2Y./� =�%es[I� P�1e�G�G7K)�nx�~�
��ۗw%��. �Ā-﫽�˜��\���S��8ŏP:N�3��}�p����r�� ڥ��`�="�дefa,��F�"V�=;{����-�i����.���c\�^�9�Z�����Z��/���oU|�6�p��`���r8�p���r,F"��5Ɗ����z�	����)�X1+�C&��8w.�Zy�L}��Rx_p���f��N�������P��U�B �`$?�����D�B�{�[��uK(��^(=/�Q�M���y'�8K�2[�EIb�g��d���,WYlj������1�a`���z0c4��H�DK�l^D�0lm5�@ѫsD�V;zO�������Ҡ�Yj}ڶ�{_���ęt�`� �^�,b��oL.x�AB�ݷ꽖1�����\<qT��:�X�d�"l�v�`�E�'��[��z�%�����-?Tf��{���s7"L��ō&���LĮ���'�7�tF�j)�A��vĀ&t��K��H@�q�@WnR��N�_1�k���~I}ӻ�l�� l��rxuط�z�RnjtB
Wj�&b5��:�Hr����]̚�#�&�E��Ke��@,�1r/C��k2Qރ����s��S2��y���(�\���?O���'yRh �!Fl������q���ش�Ad?]�+zUԻ%����5J裕)�ѫ ->���آAyҋ����Wb�����2�w(a?|�֪�U#`P� �o(��Nl� �	C��OOV��� &>]�܎~�T����}9���K}�R�S��vX膌���-�u_Y�������iv�Z��	����/���d��X���G!ޏ�?õj��� U���ڶ��E�C���w��Zݖ��A���vb�Ag����K/F�ˤ\�s�+���%Z��}H:�M��X��ZY\j����ɥ �vƊ'�( �?AD��+��Z���V�k����SL����������GW�{��
ب�Yߵ5<a�9]Be���EmWLSKT
�b�!�Z�f1��j���-Hg�r�9Ѝ�%���u2�w�Z$4O�J)Z�[3t9,�/��h��(8i�WxV��T��V,lǎ��'�A1`g�H�4�Q;��m6V���-b�8-�Y�0�m{5PADE��#qg�:������(%�"+j� AE���|�:z+���=n�ˌP�7����ɽ���sM*:� >�_�!վ�E��^8��t����u+��2��ߩ����۴��L�@�X~��M6Sp�`N�Hz��b��E��Op_z�.7*L��<�(�^!���X��q�R��
$v|31v�r�`�aU��E� ��Z8�!z������-+�׹��i>���VrN��8q4�W��T9�}���Hn��;E�7�GCG�� ��m�/ݯ��^E}���M�N��9!�4��T�/Y�e��9�ql��(�y��\~k�S���}E�����gթ=������M��ϙ՜�~"�(# �ev/|lEو>*"@Wr��_��𻧠R~D̪]Ǭ��c�����JD�.y�{wDfس��I;�]Rmޑ���P�%�m�0���&�Je���Kq �72�������f����0"�n�\ũũ���nk�o�F�Н�+���QW��Z*h�F>^0\B�C��6J��Ģ�)%���_}�Y�٢�Ѭo�ܡ�e��9T��r��
[�kG�}e����M�y/R���,�\[�v-Ga�R��I��5�S��ٙ�0�J�h[dӇO�.�|!�}̸�W���"x`��p3Rŕf*��>G� �ޙQܼ\������Ҍ�Nm���Z����G�.G�}���x%��	����]�)Nc%�M��z�03����J�w~?3Ъ�,o�~�̪�)��v�ͺ���S���Nd��W7.��2�L0�[�.�bЪ���b�?��āp��r3C�c�#[�S����#�o�5�`��b^�����%ÝD� ��6p��Z�g��ų)�Q̀�����ZϝO��>H*C[��;��> :%�x|e��HK�e�i���:� ?̢ϩ��,�}�J��-"������%���TȂ\�ͱQ؋G�&�� fz�ͺ�ýN�nNc.���X̳�R��tB��i�������?
Y0����6M��2\>��<��{Nk| 	R��*b�9���gͭ�e����HԕȄ���r�+��p|ː���y$'�詀�/z�v���Ջ�Ҍ�ڻ��u�y�2���UO|��ABm��Ū��ܗ��O7pGo�QajD
LB��D_(/4��VuJF���K������5Iv��P��0Dƺi�T8HSKB�a��)�ظ���2)]�	���]�;�^��ۿ�a]�y���gu�ŷ3|	,�sFeR��\gs�����6�+�V�v;���k���0XZ�0�j^���R��?ھ@I��W��QYʗ�w'%��Iw��Pz�o%��E�d6���*��/��|�ZON+L�i�{�tꜥ����CV���
�х�r�K�J`��}�7
N�Ѕ���6w�B,q4@�(��H�_:��5tr�e�ά��j� �a�A3�Zj� F��Dl��+ ���H4�@5�B��E�hIj�u]��ϕ�� W�� �;����5曰kMJ��?SPhsc�׾������0nį[捁=yr1!$��N��ul��N9�²�W�&b�lw���{�I�t��>Ct� �0���ī��6F@!j���%�.S��A��\e�/"�倕	���g��e����)�h;S�m
+����L�'��+Xo6D:�`�c_}��F@��<�b��1TAFsn*��[�z#�z~x�;�)��⍭����]#��K��֩e�ǎ���P�Ds�^>��S^�Zo/�����o5G^`��׼+������I����e��q\!_��F��S�* '�Bh�pZ�Z�{{
k�'�5.���TA�V�WH�	��F~2י��$�OI���%i_���Ĵ�N!1�(Z�mbL��S���f`�������(ɳkܔN�%nV[F�E�F�aI�9��MT��K�ћ��\)P���d(auE}��F�欙�W �c��K�+[o�Ф-���sq�"gy ���ǐ8f��}��>%���7�����m�����PX�9w��WF_c �E𐆸|�t٪���W=hi�D���8�� !��_Z3��-	�/��l�Hpǔ���{E��pm=���>�roթ(l���xs@Zk�w�+����+�m	eZ�²���7+s���`���l�x���Ǫ
WF�/l�6���Z�)��끾������B�7�V)זA�3o�bI�����>a��y�__<F�������!cv�X���;4��:`-�
��U�X�W,J�������.]�-^D�6ܸ0�6�B	>U�ٞ:� ��#�+4��`�!����N"���6i�t�Ӣ2_�EtZ�Q����|ݔ_5^<t����ɡ�lKK^��ݟ��ǻ���p=��q��	��4�J�SW�m����7bh�)##c%���Fl[n;	fO8�&��!ιK��%�	�ڙ��Ҏ�i�
������[5lU.�X܂�<�FB��T�!z�z����ŵ�A-�r#�eo煛��J��j��eN�${H����b��v=/��a��X+�F�p���$C)J�#U�f���M�MИr5�۱���V���oU-~��Qy�e��k���BY���jS"q�%O�0��Q�>8F}K��ϗ#W�p��6ٷ�qf\p;+�q{f��߲-�z�F��%����6N
�b=���������E�N� �K��hQR	ӳ���l$����ib��5�.��_5yx��������pcT�yY	Kc��l���M/����$u�%�L��(�d�^d˧��s?�"�#O< ��&�zAI�V��w�/wps{Α���.��
e�6 ��l��_\7���",��A����4��_�Y�`��c��� }�JX��{s��1�U�i�B��O˶��J�	?Z=2bϊ/߫o'����`�p���LN%�ی�b��{hH����a�����'�oi����2�:�YР �
��Z�"תIblH0�a�g��(v�mȊC����E:�d��J����w������~ZWp�7<��=#�����[��8��r0(ҧ/@����D{p�l�jZ>�'���{<��
}��{/��M]%�B��,.��D#�o$GtV����'��с�u�diS�#Q�٣�̸7�p4��IB�6Aܐ�)��eg���"#�l�]f���<�\�E>d�$��Z����(xcW��D��/��'�Ic���D�TT��.ʈ��wW�-��=s\���'����P`z�P �P��r5hӏAQi�Ku %� 7�f�Nŕ�WQ�(��.g��g��*|"��w+���9�X�P�I���:�.���}�{��՜���B�@u�[ʁ�p���b��>YI�~��_��������r�R[%�)RF��k��$f�f`5R{�碢pZ�>��_�'�k�+mzM�WF�Jמ�TGǿ:�]�U	r
G�J�F5=kL�9<����G��=�(���f1v��~�A��)ib$TV����>���ļ��F�e���6G�s�|ޘ`�f��Fz�=���{{���Ji�N��d�:�A�L�M��o*�0��n[`:�s#`$rWL��J`g0��;���I�;%�6v.���?��c�?����v�^�-d�V�x�wc�����[��"��z�S�v�j�5@�.5W�Nץ��&�n�uu%t�\e��&�:O�i�2|�?)a�q4P�*/�d����MD�|VְT�_���ȓRF���-.&���Sn�Iť�S7~/����VCx瘘b��}�0���[�s���a�I�'S&@^���L��	�`\�*��h�7V��-�Y[^���V�l���D���4�����̏��f��QT��_����t���t@�b�UҹZ�> K�7@Ķ�?Έբ�����*�õI��-�
;jơu�/ٮ$^�5'Y�4��,��cl���ѩA��#���~'\
*�v�g�J�gZ��kDu�]��qo1ֶ�����$�b�ADX���	��)�/�٥�m�z�ùr*��$񁀕���13
��Ӥ�B�pU8��e���P�{�-��]��`G������������VF���(��m
��ȯ�%BcX�d��8$���R�fB��xC�IĚE�
=W ��AF�@�l�^���}�⊗cu&�!x���n,#���	�vII%Li�����W���a�����ׇ!D�����uR��{mn���pM����p��.�,{�����6�I���yaY�놅k�&$Q��x�>hC�+�a �,;J��2`����Y�r�&$}��P���>Kcx{��+)�x]PdK��xix :T�z:�%��I�u�N��-*���vG)`��6t����0�X�O��Ӌa6Y�x�];���|��GE�&v���7l~�A�r��8'���f���;!Y����.�֊����b�H>��I �e�7��t���(I�DWodǳ9X���Q'Jp��;J�������H�BwԾx�
Z���}=�s�ME�AL��B.�{���Uw��YcP;�3�j)�)�����Oa�^bMJ�[P`��m��J�k:����U9��\���4�"�A; ���k�8\I��r|����g��)@�[9�z��7�Fj���%ee���N���;��Q�e=��md�:���*Ӹ���0�nP�c�>qc��~털��>WZ�"�ymW=�M��Fy�ŔS�>T��O~H�kz-r q�B�����	N2�.G��̻f�3�)/a��c�ŭSxH�G�z�`�Z���o%,�=������p¨-1e�Q��K���W��%�DH��J�U-��� �L�Œ�3Y��+�O찌��#����΃���o�e�gX�J����*�7}����ݮ`��C@�]i�� D��(�����t�e�S�T ���J��Ϧ{I>=,��U� �$�F��62��j^#�+~�,�s!���컼�<�)܁�% a��"�G�-��w)�(VrWµ8z�:�-�E�E��ņ��|aQwl�eX�=�n�ή���Q����7����J��z�<��q�8�� s���6'�e���
g���4g'��47��yz	���v{K`A�L{�;+̐����S���xPc���~�V!ꕇ]A�k�d9��hy���./�hDug(r9�"9'b�.zvچ�l2��t�=T���/p��d�Ź`ᙓ��7[*2G�X +�����=�ʹ/�7E�dr�(�\#^+>b�q�Y=�@LF�5��� ��߹���:?�X�3��{�򯽬2]W�T;r��&L�:�'D��!p�9�gz�r��!g:F�ؠ�1��x�F��s��;�/�3:�^���5�z��@;c� ɓ*0����� O�}r���e�,x�j
���\���_A���'��{��ZXP��6�Z�x��.p�D1yԦn�,��zL��k��z�1.���Z;��{���r�A��p�X�ǥ��*I�n$p﷦�HmLJ҆*��8����R���S��i/`����E`�����h(0����i��So���zh%�����(����4Hz̬ǭ���!��e7\�2�y+�f:#z�^�����K�:����|�mC�DɏA}P������{r��``��px|�x��\�伉^��eoN#��).�M���:�&�'j9����򬯵�|�*Z�ն�Z��K�w��z���Su�Ez��A�@n�� M��E�jTOh/�+Hl�-�-�L̖�����?CNmɊ����}Q�@�4#�s�i=�'t��7.��^Ԫ*6�$�)�q(ќ ���cK5R[n��X��w<�y*�D��{��c���N��@D�Η '$?��5�A��S��n6��R��o�����M򄵬�p��/5��[3p�Oj{"݇"�Q�����
���6v�Q0T� �8$�Rr�͡+��bHK{ڜ�?q<~w��^�'��8�L�`:�>+(
��z��ӈ�w�j�3R;�N��H]8f���pb�|���"og؉�4�fe��|��[�(
>�I'%B�F�~��l��[�:�ڑ�!h9��UD���DԌ���RE,G��i���o�hq�i��3���[۠HF�i9w%M��9�{w��=��_I예Fw����X�5�7���,H�Q�OF��W5M��pL��n�o6I�0wW�*��� ��AS�ro�W2(�:���c:Y�"O����5J6�6΍���TTY��'��[��9��i�
�Y!��P�{�L#gP�_�1(�G�G)�`� oM��F6�y��K����C�۰Kua��D�����3���M%:`f�P��/U���X��hS�
5�U��KOZ>O֤��D�ha66�f�����~�Z�����7�tK��(в�&|�͵�	�a^�<y��L�^rԮG��S����ޣ����Z1�@|��Kq�a�Q��S<��)�^�0�326/���q��=�R����m\���t�Mgg��+B���J3  �(ǥx�ŋuW�R�M� W��i�8 7&�ƩN���Sz�
��"XZ:~�8�1��T����v�ړ�OpC�2�h+��fm	q�DD���ڄ^b|9��g3���+�L��b�Ȯ�۔&���-&֓��!3>n��f���I�o�R���e5�� ��S��%��I"�5(-O��dX�Q�Ub�hX^ 40E���҅������������:H�k��J沶���F�5�P�f���v��-k9f���e��"�GIm����QM��ފ���So`����'��Y�cT��
L7_ݑ�.c5��3#��u)��$�o��)��y[Z��d3�b�"���^K��+5�DU�s��5��fⶠ���7Q]��hJ�O��ߧ��tH��H
ՐR�r��FqPuP����|�Q�*vAQuR�1 � V�����r���źɍ�Tm���� ��,j�5�����P񪩽�h�&/?|޿��{��܊;���2P�H8���f��>���%ӕ5Gd����Y4�iEo�ܒ��o�����[O��/}+V�1>\�mC���������ĺ�yp��B�S2���42d3&������r���*��_R���\	�'U+?y��x���s���2���|���s6!9�䘁�x(ټ�o���T3Y�{��,}l��4z�P�W �#� �'���#��/���6��z��G�nO5�M�2�($�Ɏ��M���E������`:~���*�3L��"�m��}��D1p�pW���,+�V�v��v�&����+QT�&��j��'|O\��^�6!���L^��D����w!6�DkmA`�_�Ϙױᙥ��������ք�5%�����nhli��j3�fߝ@Z�q��LH��?�LY�/���H�����]q�.����80��D�A���HQyM//�K�� ��ꂜ�!#���P+ɀmK6"��¸��k�q/ʈ_��tϽ(�G � �m�e�����T�uh�gyQ��k�ϓ�����:���{�-{Y#���x��d���Mb 5���N視���E
]Sd�j�}kpJ	[Z���/� 6v�ѩ�9��� ����Z��'t+�p����w��A߼Y��J�-�4R�:Bg<�o~.>} v��MD@�4P���6�گj�ηrk�A�A�-ž^�4�B,�R�+�@{^�Ƌ3�~�u�މb�#L [�v��&���9 8ye�z�ۇ��	)�L�h]l�D�Ay����������ܢ(�a��F�j��έ$�w�'.w�D�sQ+c�M�7��j%Y�8�� IU��p���u�'�k��i����M��gV ٚ�Er7�^����,��8J�����U9!�C�5�u��~)[���W�L٨«�z�8!����T���v�X/d�Cp�B�2��(fg��Cd�YK��̇���#3�s��A[2��������G��ZR1u	`�^m"X���j�:���t"��wA&p���snN� ��M7�c�u|Ʌ`�
����K�[MY�g!�St'@k�u4�@�d���}����&�]b��b\Y��/�d�߼*I�2������	�I%WR6��B<�[��]�G	�����MxJ�{\���ld�������YO��G�?E������KA4vx�i��^_�z��F�����[+�ᠾd�FSf�U�9��u3DKi{F?�d@ߚƐ�g�;�E���
	����,�����A�J���q��㿗Ԃ:b}���s��ntKbE���=�͏�TM�#Z�X8q��`)�ĲO���S��á����
���q�{���3��JF)��)pI��M�˴A�4�}�`n���
����E�l�).d�h�V��>h뱽���Az[� ������L����WM=���;7��M�'��VN�Ц�Bi�3�B|
�C��9|��qv1�`���t��ɢ\��+ΐ�e!۸���G��T����}.�hi��2��-n�V����2��h��f 1�����'0j����7�,{�����g���R�(Ӷ����o�3K�16 ��y���NJ3Ɵv�v��c�í�5,��4f�0TL#s�;�O�� ��ĭD{Sల���/o�b�\;��� l���KG=wcR�����_��W�QN�	�)���%j�_ ��@�S譛�-�yQ�&2���𠦌��_}����|^��|�P��A
�kS��d���d}C*���8�|TD����ֆ���[��|7*S(x�?ͳ7 An��������Hv$�Y3-ܝ{oP.K��V���	h!v��$)n�X���$���2Z[_Ԓ/`�;KO�u�7%�N38J����nm������+��Ϭ>���p�����a����L�5�J�z�Q���dl7�QI��:�oO��YC�
���c����D����� �	xb�&�1ED���J��T�3!����'��屴��Y�yq��\Hw�V���>j�<�Q����{*:��了�G8@c��p��/���"���J3-8]E��tׁ#,�U�V���J���IJ�]�j��������ֈ��?g�H��
����Q�A�H��˓�r>Yn�k�D��Sn4��|�
>=���gQ���q�$�*T%�3��s���3~S�k�F��U/��WބCD�I�������1��P[��c�=��Ǻ���	��!x�`�8m����Sr�Y?n�d  �w}nՆ�L��F����IАNж̻�"�ɪ���w�9�� ��(��G~=�Y
F7�� ���\�h����3��z*!�~������=����oY[fc������e��Q�wi}ߊ��e�cۣr>	�Gg(S��ܖ�=	J����}���x��D�hVu�a?�#�<q�-2l+��� 9h�4b�ӛ`��!39&�
5�oT�� '�B��G
5��F��wv5 �^U4V�y��in�����Еo��A�'��%�l����<���>�{ ��� [|]ޅ))n賤���\��������%���)$�L�c�Q}�F�u�(�.y�7��f/ٱ��q+��2%w���gK�R�����rpjU9tE�L2�Gc6�.1��#ɴ������� ���#b�<Y�Κ�c���c���X|]���d]i����Hw��ě)����w�F��!�����4�_��e�ehOO���N�(���i>�iA��C�4��6���*h�@�=���q�oDS������bR�����G�#�-[�;e`�ih&���=4���,���^�=MH|\/�7��U_�Ư)D�M)?��$�ѹ���1?u>��Pw`rAڸA����}�KBe)Q�k���
Š��S�ܛ������/n����c�	=9ِ�:6t����9�W5�%R�j9=I�N�K�'����6u�Of6�L`땤з��P'~H`�8�AL�
�a /�C8��E��� x�DxGen,�H�㳉]M�/��ga�5���@Wnu�ida8���;���/|0�;�4�m�u���g��+�˅a8�F�Hˀ�0Š�7Cs��<�0"��R��0N�C����~/�nI�/c�8�_qZ_:�o_SQ�V��yۗ�A<`�>t֠���M�IEc��/T������'�9n</l�<���7ȣ���=w�S��uI?n� `:����9�n��<�;i\?_�rr^�.OlS��%��ՀK��Fm��t��=�ͅd%IS�l�bX������廣���&#��ֻ��lb�(�w# �X��D@ך���g�����Vyf��=6��5����=�zq�t���]_��^r��f���zt��ގn	�^�,RD�*�_]�uҀ�N��c�Uh�|�ՆG8 �k��*�27�s��~s���/Rٜa�bAx����Q�{NLU����B�~1�(چnK�){Fk�zP��7s�8�;~���́S��Q=������ܜ?��X���_������S\)C4�������8U�dۨ�[#Gq?�>�����,�N)��2ZY�=���ϋ�A_`���f��"Aw�3���V!z��jq����v{��K5��`�-� ��sB���2UP�M0Z,�G^�m`���4
I~��SI�7_9J�e3�g9щi_ �tв������ڻ���A�?��H�xN,Vd	!���}���G�Fl��8\`�U렳|c�9�唐5�eVn"�I�����uW�ߩn�O`!��
�d�`+ؒRPKks�m((�3�GI]RY�mЅ��v %
�U�BVZl�|�?�|<gWɸdu�&� �!g���6��X��
0L���?�FR�!t��&d��?�K�ćC���f<B�r�vM���43����?��]ٺ�d�2ꀩ��;k���9�1i����S �g�o��[2iW�:vb�		�����a:��C���*�BN~�r�'VH)�%�uk�(S�%�m�B�Cؔ4�;��~���J�9�kVLMn�izNa{��OZ�#���p���H��̥}�œ�7�4i�����A�f�cp顭|ޤ�f5���*��R��|O��-��^J�[����}�đ.>[�XRi�4�%�d�=1��w�4z5��%�@D,-<�[�4�4�r���v�lr��>L �|��12;b��y�Yo�,�(����SA����d6����_])�R�[���4��E��
U���Ҟ�#��L�{���󥖆`K��@K�Н�����ZB"H9_��[k�W���@P���M�W'�l@���Иg,O�1Ą�a̿���V�洽a��ݧ7�����Z�8Y�M`s�71ʗxG�=wb�y϶}�;��=9w�>�nk�Nt'k��K rNv��@�!aZ��f�3�lw��Y��?������r[�N:AQ]��������ʥ����%���T$G�̃�M�$4+�u�- ����|���n%��p��D�	��'7;�������ǵ#Y$�r�cd��%�d*��e�u�*�
"d���N��&����y}}y�j�N�WC�f��%݄�;���Ɵ t��G��SH�f����ktj>��d[k�e. ǧ����4L��=(��qHv�^��A����sl��(��/1������/���|e;,��$��3
�~\�%a���+E8�Ó����q�H��ڢ�1\X-K�� ��J5�3,4f\��;��,�*o
��^|�~E�S���ЪJ�uVj/*��V�W���,�g�m:+TCE����G�e��!�U���O�NvS���N�`7����-�J>l��SQ�+؆���:��k�����	sf�e*� �r��G/kc�s���L����$j����'�����C|�]��|B�(�H� k%��J�/��E��£��.)$�o�!�v��[>�����bsW;cL�1Į��A	���.������x�O���<S)��M�+�J�uPS�t=;�31�fH��b���㭚��bpHq�
aO%W�|��E/I��M}x��&5�#��:�,�S�V>:����$�J�z����	:9���Ң�mS������T��͛���~�q�5�9��",� w��[5�z�#��T@T�[C0�l��D�Y;��`YAZ�b��6Lj�7^�6 *��C��s\�*O��#��g��I��@�
w=`�r~�����Z�93@���7~/��$<�8W�q;�t�
N�k�]�alĚ��+:ش&s��$5�_�k��Q�����u�"�_�ڋ�	���he�q���k�B��	����1�4�_�y����6��/b�[�J)�<B�V.U�6���EZ�>C��/�ղ67&�s#:�l΍&(w���S#�g7��CG`����iW�c���sO�ox�
�D��M����f�ѱ:jy�:�ޔ.{ ������;��,�v�� Y�w��`�m����k����=�N_�J
��#ɣ�Z%�b��k��xr	O�Z�ǐ>|}vi�H51iV�t�3#�vlu�8��l�� �V�f�d�[�H6@UrE�'�tb��3t�ҥ���X�9�a�!%8Ia1�9���-_��e�7tRd\����5�rE>�U�?O����D�`���1�Z���[~h15)�}�C(7+8{FtZ�k�:E����_�~��9�,�M&Ҥ��}F���!�����j�����u#*e-U�o��ג�G���?;ޛ�F���~���#O>b����Òh��m�WK����@�$���⵺���?�`nl���wr���@�l󻩋����h-T��O�X'�.�q	�<��$$)�}'��p�[f�Eh:��Ln��>w����p~nl����^o�:�O�
�N�#����.+ص]�e��Ɋ����}�&H�S&�%�J��5҂iD��>�u�Z��������H�>D#D��i�䶱��
&ڪ����2,�$�!��W?ݢK����/��Τ�uI͵3�Ć���@�M~L_Nm�x ?o��ӧqG%G������n���ךʋ��d �M�s�?��&�����z�zJ"�0�z���K�m�ٕ���$j��qVb��I�f�a�(b�q�R P��� �����Vj�����![S�|�3�k�AL,c��� E<�T��@�5CA<�i뷐����{��o0���imΗw#Z���V��s12���!B�d��$p�_�v�� ?�EG�������f��	���1O8��@�Y�~��O���� ����-A��@8>��t������̶���*4PHm�3�v����Im@�v��~�d���B������8l�A��T�Uw��ퟆ �����쫜��l4C��01�/!����F>�c�z��I�l��lqQ�ͰA�����lS�+����t,.^ �Ю}�R��KHfJ��Q�R,��<ЖF�_��\)�e�a�~�I��d1�'��J�W��d�p+DE�����q-�)ٍe����̵���7u]o��ʥD���p��$���ZtU������C3`��)mF=���n�4ԑn(JG�[#<�b��P"��$��"7
nc��X��������5F\3���U�q��T�Mnk@RKD���}����%(x�����R�^�.�y��{��$;ơܒr� 2t�_��szِ�d~i�Y���/3݆���i����k`|�2���	��;77�=�� �.�w@m�!�p���x�1��S� �ukWU0j�*թ>5�oOa���}MƸi�#[��!`�G:���DD�9υG�Rtb���b� ��;����)��w�a�{	P���������ޏw^���2F�`Nɒ}e��8m�Y���3�iW�hb�6:�oF��pOI��< !���ɥ�F${q�`�ŷZ��j[�s���צ�t�A��_^]?}*-�>L�i�0l4$U�U��hH�ݼ�l6<�j$���
|d�$���r����ңX�\��$�$����YEI1��<	�"b� z*5���RoY�-4K���g5���gF����aץ'������<����|�>����%���'h@+}�-��y�h�?@cvu5�zx�p�!Ɣ�J��4�Q�����А9kf�>�W����|\L��#i��J�`�(wtb�m�" �Ǽ�
5@Y����˶�amf�˃zao�UK��6&q�!�6�mR�#=OW��g���c�qh]fn�v?�M�����r0��h�8�;oO����,JU4�� �I�L�2��%��A��-�}�u��,g�!�(��Eh� ��?��4�Ȑ��gx��� ����s8n�v�V�?��w_$G�+�_��b�G��}$�_��X�t�i�t2���x�qa���(ʊ�L��kuwM��BMg=��0���ā2	�`�}F��m��B&�Ď��j�b�<m��-]�^�����J&O����Ǔ�A_�3�V��C.��L����@�p0-,�}�c�5ރ6n���@=�56�b���<"h�Xҽ�o0y<�0}��g���E�oRBЛ-#�O��QH�� !�,AF��'oA�)��zJǆ��㊙������FU�� mVS\���+G�f��H�Q�w�BE�]H����|<�_����'�P � $B��G����ݰ�{c8���Ɩ�8F3�~�bu?P!."4v�%���GK�wm���R0��O�%n�ڝ���b���b��₤��f��ҫ�!ٱ�{5���f2�[i��rj�,s!���B+�/�ɇW�#��rW�1�l�Ȕ�/�>�v��d��L�W����
/P٧��۫��d�OֹЎ���"�-b��S3��p�6@F�'2�������7�G�y �jHő��D�֎4����w9��g�༅����r ]aT��æ\�[4�S�C���M'h=��B��\��0#���=3w�q��4�H�����,�e�C��q��YqY9&DL�� XI� `�3Xh��!��	ӽ��ў+vu�٤1	��{�,��7Ѵ�?���r ��=O�J�\��I=\F�Ou�� o�J�<f��%������{x�璉�9`�}�����.�̊8@�\*��'ߥ0"wFŁT�$9<�訅��`�yc1-��-���d���۴U�Z�ɛ�"�A���F���@����pb��ξ0��'Ħ�Qs6����q����ԤzL�-�����xbE�n�SqXـ����Lw�6���A3`����.�ZcԠ�S�қ�.�ih�T����|�u�� 83�RҒh���ID�� =���wM_->ފ�K��e�MF� ��N�Y[瀕��S1s��h/L�Vo�҆������t�I��u�i�����>'�=���'��8�j(L #TBh���t�Ɇt���7�cd���%�**�b�gb�qأ$����*��L���RP3���]�#� 8� `�d��(���s�(�&3��������VUؗxy������Q�T�q�D�#�M��:~�*}���m���eIm��Xp`v>)Q�tU$�<�dt�o�Nف/�ҋ^X.$||-��縖1�����хd"z��8��3�W�z�i �xc�\��^��k	��K�����[-��k���K.��#Lg���jC�j��8s��z|�a �����Ņ��Wf��mHqku�2�A�,���},6�=��	��٨��^q�f���k|Y���-�lU^NU�DaA�>F��J�H,ɞُ�߶��%'���x��GD��Ӯ�2W1��:��z~���E��k$�o��:�$s�W�I�>��(�ŧ�OL;�{���q[g5�'X�R�p3[WZ�`�	K�k]g;7��`׬/5�%����Z�׃�@������&e�4�i���\��Z�X��ڶ�:�&�����aN���@e�3zN�V�������Ȱ���?��)JQ������ �$�_PIp�9~u���
W����M��mnE���|����p��;'mD�N��˿�����4�H�m7r���9�f��,��FQ����z� �1q����㠿W�{�Ȁ�!.��|,|�y����+�Z�U"�X:�?�����M��ո�ɵ�lGʐ4'���B���G")H�'zP��'	d�ә����;2��]��?�h����Y͐��/졒"���Ij����f)�/�B=�:;(�k�p�f���?KĎ�Y����-����p��r{���<y.vn$Z��3rU��+����+W4r3�?�뇯�Ca�þIm��Ť����͢���D�u��0~�F��[�B}S@�?���QvwJ�,��?)SAdh'��Aa������O�/��,]v�Nc(a�E�5Y>�]��Fn^?H���8u�����=&ye���a��(*�=Mv��p��Yk�����i�R9O�{zIp��Cb��z�ּ ���w�ލ����b2��E��� �*�:$��Ȯ`eQ�8T2�Ea!��1�e�.���a��7���|J�v#hK�w��R>7YW��"�f?���V@4�� D��J���}r�3 O&��-��,�!->-e̳��k��PD��L�F������^��Pn�cJ��ȳT�v�bL39y@;��`�0�Z�)��Ѵ�מ� �\�apD+� �P�xZ`�H��c6��X&�ŝc�	T�)Y�3�Z��Ӊ�����P���Rj�΢��@QF�4��(���7؜0�~]|���c�Z��d�9=�d��*f[�4j3VD��{>!W��ƶp�.�n�(vI`��F��E߮��?$W��g��S�ϖqȳ�KV��ω۪v����W3Z�5p�B\曇��{�t;�Z��5z�o�h]�$�::d����5PH��f�*�����&����_lT��aK��;���L����ZS�((�0�m�U�����E�|(���3���9��G(�������{���I�A��»��Q��aZ3��]4p�Z��F��P�Z�Cў���.T+7�"T���/ȃ�״�U�����6��r�y���l�gQw���e8"F��@���&����s��5�^5E Li��k�a�g��h��mVb98tXӏ$��z_O��q����Zny�\a;�&s���묙�nt!�\�ǏN�~e{3Mc�W��q�\����mT���	?(�}��O��QB�Y�.(�		�t\(@r���N�i�<Z�_a/�d�G�u�g3xߏ�&�y��F�|"sl�0%G,{
Q��3���9p=CnB�j��u	@� iN�&U��\��7c�*�p\"�郈|+r*��ka�{rv�<�z������Qv���d"�H��5�hˇ�ЎM<ţ�綱��HA�K$����q$~k��<q��aF����r��&:HÂ���cǋ���H�B�06��������Α�j�s��ѳP9�:Q3��Ha���+9_S�
Lu��{bSdy.��Q��q*[Lk��=��p��.�-�^uK"s٢_Id�!XQ��.�z����+P�|&�0���K_��1_$_�	9 1�Gl*K)�F�?��+��u���t��խ�N�v����t�n��Y"G�f��q[�/Q>��M����]eθHzDo>��U��m�_�>�;�o���UYX*Qз�:GŶ�$Bc?�]� �r���С&�4����*�:��`+lB��OO�o��9���MK��#m	��	�ߋ#����%� :;�� �5���X|����]I�BzA��>z�nQ�6�Av\vM���-j�1�ԛ����3��PI�j�.�oi�B}y�3$M5I'����O~�W3@�S�IQ'�I��L��7F�' |{O���'����A/�����}]�Պ 2B��K�����PJ�(]��Q�`5����72R��(�6 �5�'�S��+a��X�}) �J��(�92���{�R��'oz���AU@���N��bk?��;���n{3��:!9��V��ty��G[4��}�"��J*��w¤����|����b�M���� j�4��Wk��B�4�)������q6T���j�~X`w���VR�#�k�hG.P���W�!��j7��9f��?�M{@I�U���m���j��(l�9�7�tq�O.��;�6S�	p2���@b�v��|��㏼�H�������mx���fX��S[b�`��5l��N݄��BS�fO3��ͅ�#@Ƅ��]��m����a\}�U��/& ��Z��r����lɔ�抃b�>F)����"��#^e�p�

��篟Slȉ7��~L�ub��ב���m�9c�F�]%��3Q�s���ˉbLV?�0��A[Ix���u~�t�?/^�$^d��+�5G��q�$!9�B'�d�(�8rSb^��+�����T��_��gӋ�y�}����@���	}�j�_$g1�Dθ�/�G�kU�BB�1�M�\�t�\7��^���Ĩow�}��h2�{p�o{�6='+
�o�qo���C�4��K�m{�Jlu��R@�D^�dӍԇs�0A�E�t0|.{!ZA�OG&���TA�?I�MO[�g��F}v2��Ky֩iK�f�ށ�����&[7e�(�8 d  s��;T̢u�Ή�epm�mF�X�Ȅ�\ ���9�Θ�>υ&Tt�K-�Չ�D�o�H�Z�$7��V�+�Feڇ�Y�������m���Џ2�A�fDU��F�4�φk�]�G]3(�a��{�UmҚ���`�3ke<��:Ѡ��ӻJ�������i��x�ܚ6	D��1u���0������T�
댬M9�LwR�{���1��s#D=���dG<���2}#3��4�5ϔL�5&���VpŽ�8	�5_�:Re����u�Ao�	��ٵǚ-�KK&�}e����)z *"S,\#�J �k�PD����Xw�A��#��Q�a�$-;�Ka�&��D9}Ei�Ӵ��7yTk�#X:l�ҟ��nˬȣd��w�2�]N�yy�V�$8�0���;I׶��}qM3jJT���Pͻi���{������G�ߟ&�pb��-m��j��g��\��`�x7pX�x]���Y_Ur������'A�������Y�y�J\ߪf����!�)�MoéE�p�3M�G62��OvI-V�����tݐ��4W���B�Y�x��_z��7 à�L}HJ�<�m|<^gۦ˔o#�F�H�0F��$3@��>�5Wo�W.`���4X��]�G��\Xb���dw�ҟ�Pj�]$���Wȹ����Ԇ����Q��!n��NBU�!����];��7�x�~�!Fn��CeM K�]��vh:��I7�[�f��D�l�=n���%,���Ւʈ"ǫ�l����!���8�������H�3K���W.�����I�]�Scǂ��s�<�F+��Ǹ����@�I��}��;mh;��nn�q Ek
s���-0z�i={�$B2>�KL���S��� h||,a���R���.��7Z�$�1+��W�/�ט(�9�6�I_�VP�9�"��e�Bizjۮ#j�A���]_�im�V{�"S������;�ѳ
�@��DOU��>�Z�5!@� @��5�ER�J�iFG�#�^zB��������XXr� �(��Lc�d�~��;U��S�&���]�Ū���xZ2|i�j؅|g�si��NA�=E.7C?$\��[���sތ������� ��P�~���C'ʀ�3��w6-#\E�3�%��=�I\���o�٣H�Y�/p�='U��h��l�~=�+�7ni�L�g�䚘���k���~E�?�~���7�`f�3j��ě�)� #xB�uO^�ң��H����N�����`�����!����ɛ�B.���b��e��Lx���t<�Bfdy��|�nl�N�%L̉����d�W2��
BJT��b��h��f�D�.���0��<�,WJ���Z{�+`$��Ps���)s	����Ԥ�����o�1���y��0q��Y������v�< ��o��+_c�9I�r�f�|g�b��PJ-�U[��p�t�����{z��@�	@=*��DKX���2���0Ī\I=��-?=#���ne�qf�=v�L�%�����N�W�ٳ�Yȓq�붪���F�FX���6�ĸ|@�&�S��G+��7)�kU�,�~	�hۢ0 �+z��'A�D�r�,�LȚQS���H[���[;�m¢�`���&�&�o�)�
�g�erm��*�����C�e�YA�7�$�Y/�2	2�4�aq�~�iw�H�Ypb'$3C+M�F�]�LaTei;�7#Ŏ���ҕ�2������ '5j��U!0����JHXu�%m�o^>4�K��'j}G��'�n�Z��E��6���[���O���Z�N#�.���Q����m���.؀���l)����6������:�A 1 �b�����@�2y���ڮ<�D0�q���đ���el�t��Kt��b�d�r3�I���*fqw}�%�t������72�K��.;�q73TV�whzT�*[ �x~؇�7�W�l�]�`x/����F�C��),����ofr)%,����1���x0%?�q��V��ʁ�o%;�f"�a���`t�-��g��;)�O"@��p��D)��Q?6"`�R,Q�ج�$�ّ���`ZS��^R�FH��!�\�̀�aSz�� �ن�"xhI�	>
�@B6HV<���Qv�]��>AQȸ��"�n��o�w��E�0Y]o�p����Kw�K'��*Sp�t�T�Eag�a�=�t���ڕ&G!�I]�x�,��7�.6ؤ�[(�4�W���'*�z��V�	%2+��Pz��W���\�4�Q����͵�֨ю�/�b[g^
݌`M��	^b=3�p�����}�v�((�_K�2WvF����X�]����;2�RW��H�,Rj7��֘���G:އXb;E��M���/�
�J���:�8��!+/0�.��=x����"Q,Pg3S�B��;��{L��g��s�x���a�^[��$������i��a���4òE�����*y��e�#E5��wW��Z�2�bN�:��^��d�B&�sݞ.�g�E����E��φ�f�Z���	v���2f�|m�y`��2/���=���m�>{b�٫vҙ�-C|n�+<rwo4E��j�|."�2J�ߤ������{��r��yQ%E�((QR]!}����:Ô[�J�߿�!�����E=�_�D�o�!�NG&ۦ{�f���U�(����m���!��B8>g��W3Ӂ?�3S�2?̛�llm���g2n�cel�HU�wX����
�b]�> ���s�i����Uב.��ÌS�V6C|�D����ͨr���ݯԢd�����RB�
7�Ŧ���-��������'���1�ޭ�,�֧Lm
ś���h�!<!�\'�����d}}��P�_TR�Sh&���V�u�S��º�oDg;2��5r5Nkn���E�N��K	u��v���I��-y	��je�#W�O-o�Kln]X�=bQAiMS�DV������-���F)���')�w�<V�=a�/�Q��k }��6@
�W<��r�~%:���E����t��^IQ����ZB��2�W7��PS`�ub!8�5;����V&�r�W�2�i���3	��q�0�����ע���9�t�)�C[{��1�#�Xû� ���?~��F����NQ=��-�\s&�s�����?u�m:��FM��oP2�>$O�9�G�&���J�/��c���V�����#!�Ĵ��pӶ�P
A��U����V��TTu��1֓��E ��#`��,`� ���"�ԖL��%'eLq�]S��@{�]���S�a�/����O~��m��,@	u�_�3,0S��u��L��o��������$;�{O�7H!���U���<�ݰ�!6Xr��Hj��I�K�0Y���'�m_�~!ͭ�-�M\u��@�N��b�2;�-t-�p!B�u'������)I4�5�{P(�H\��q�m3��W�jO��
���HM2m(^��wUۨ�̗oPÙ<1[�p:�]�{���/� i&?�&b:�E����my����w_h�{~Pk΋;��qz�Jؐ~��Y@n��o!wQ�T�q%�w���6���Wa3AՊm?Č�o!�l�g�mI�aT��^G�d��'n���v���:<ҟ)jR!�M��웃� �cu�28F8ϵ�w7)�2jw�����T)ڄ��M��(]�� N�i�f��y'��̀�s3(�K�%H�Q���J���#,'+�#��]Nk����"8�bx\�ccO ƅ�QI!���8z!�^�+ȓ�f�}#0�rj}�n���M	�z�R�Ŗ�siKW?���"���B�֒Ӵ�{A���ʝ�dXgM�Aq�c���ԫz��H�����x��0�Y���P�%�+-Q��
�h�t�5����t��
��(�X�U�tj�@]����z��Z6��ɺ�p�*�7eCE�M�3J}�[�O5�_hՊ˩f� �
�F#��ɀ}�!�
�<���#c�>�(��g`��A5g��9��+�c���+E?e�7wL�_���"�Y��j'�$B�C��ӟ1E�GGN��H�ȣ<�g�{Z����
�}7y���ά���\G�m�6f!����'�̛��a:����qsM�w���"�հE(�N�c�����\�O��^F7�[�����s���K�<FJ��+\o�>P�Q{I��N�#1���[��T�������w�?s��L�_�a��\OY,<�s��̱�$�kʡ��(�uq���o`���ѓ{�����g�r���z���z���)f���O�������&y� 
N�Jv�_���1����������tBME
Q@���e6��v�w�*H|����[u h/L0�B������Y�Ded��J����Qn]g[��{��7�l^�n�r��$G�>u��>�/i�}��Z;yI7_r���ȾI�i��*�\J;Ǻ�<��m�$,�fqQ�gf}�.��L�0Eـԭ���[2�T#U�rd�@��n����n!Z�Jp����%��w.�ˡ�>|�q��l��f(�}��a���l�Y�s�r�g���'$x��2���r��#ߺ%�M�ӣ�n4i/qh�
�4dw��D�^	.�^1�[Q�~��i��Fe�f�,�"��x���	��-��|�`@D��M���ف'?pH����Y��h*(I�I�6���f�d�0�0�m0̳B ��wU�)��Ƈ�'��,tK����5c���hM�d���g4v�/r�ԍ����Z <��M���n�p�.�% }_K�];�gB�߳�i2����#��)�%�:��7��w.$.�%K��ϣ6Bё4;��))EK!������0��h6|�W��\N����q)�\٤zYw�7�=z�X��_y�~�g��0V��|�7�S2���+�I~)�a���Ȥ=8���Q׆P�gM�`Y��U�]HX�vT "Dsȴ g��;�|!����zפ:���𛕴e~��c�Fs��82o�� }������ �.�DB��H~ko�Z��i�Ol7�.�zVZ�ґ5I�*�-(�!�ÿ.�^�	���<X^[�p�ϫOٲˆ��x0��N�&�4a�̄�k�G��nо�&����pւ�Ss�h���K�bE��l_��W�Ư޿���glb�,�Y|A�a%5f���pj)�i��#= �����|��'���� �r�g^��K��yE�z�b����'��Bf5���v#�����\�cփ��^7��-"1ʍ���|�zv�39:	wW�ggxr���[�O5H�]���ϼ���6|��j�qo)R���W�Ѕ ���zxY�!���<H#�����/�R�'���[q�6u�j8��Q��0��ĦϿknVߙx�b���󨘶[x٥֡]�.�U�;3K8�>����?�b�8���_�����+x�E���Z�XsG���G4͓D9���梋U����@�w����kf9O�(�jZr#���&؅3�;Ȑ��,
�������J`� �S��M�t������m���'�m}�P����-=6��2��68�`ԱAV�V�X[{7���S��k����%��A���g	�=^_>�|LK�B_7�i5�M�_d��C$�~�%3�����G��R�� ��z8�}5�l�<�F��`~�=�5q�ذ�� GiG6�@Ͷ�~J�G�Q�X�Q	*�g�+L-;�\p�~�O��p���<�ak��yJ*�i%snT�В�x���\[v�����G���#E�^#��yɆ���~E��b�WP��U�2��^��_j�����B���e�<�CCkة9�Z��ԃ��H�G�`���^�w�Plܽ0>���:�_,���$�N���ߟR��Sv����?z��g�*�X�B���]�%#�=���ke[=���k~���G�Τ��C�H�{j�F����e��F/���d�YP�P|�J���	�0�<W�����'�� ]��榐z��t�A&�����U��Nܷ��5�c�/b��#�fZ�0[�h G�R�1$ڊbf���yS����z_�DX��Rm�.�_���=�����{�d�SQ�4/����W]�{?�n���T)]�^M����Q�5�}��%t%�/��ɿ�F�oD�?���+X�D ���(̻��H恑R�ɼ�=
�������QH���3"��ȧ w��%յ�b6!�P�)�2�a|�~)�	+zD�i2��\-�l<��A8h:�Ck���?a��@���vL�0�����B#,�hk'���
��q&&�R#�#��S�g)���d� ���G��i�2-�.L����~"�sjs�a{���֓� �'�v~|�T�˼X�Ue}/�ghu���$K���� ��Qҗ��R�'3P�r^Ft�z*HS�ز�=�U"pS1�(���_�-N�
Ϯb�W�lG��/z-n�Fh��!�Y�"�1�χ�+��\��	���{���h9@�ap�����$����ì�޷����Z����̫�,*J��=�1_���7틤~ �|�ݡi%AUㇻu�4��;�S��C�S�ڼ���;i�[^@Y�Ū�����.-��ʬ]Vcg� ����l�"��*q��hb-���>���;h�pH�
[jA? {���
�f<0��8ǽ�zP ��|(�`H�<W���4X:4J�'U<��o��ܙ��7�U@ŝ`2?1�k�KN��"���ֶ���-�1^�^��|+K`>Y�$bq�(Ӊm�Hc�٘Q�_ǔߜ�]1P�!�_9��RG�"�sІ�X3kd4d;B��F�l��#�P�����)?��RӠf�eY���r<��LLX�� [5�s�DW������ݭ��ե����?=��U.��^��(��ojܖ+=�Oƛ�oȊS����!��� HX޺rɵ��'52�A*�{�%����j��;ڸ0Lm�|���F�M��/˧/4�~��(P�:�2�  �l��_V(|�p�j�漫�m�:�^��
9ߡ�c!'�|<Hyٸ,�)����2��@��� �&�ɥȃ�.�������te7I��������"2���%��S������3l��HF��\_6wk��>�]ꦌ�	��Z)�i�-��x`��.�!.xR����_�)�d9Z��*x���V�a�)�3{��AL���-�k#�3��5��}z=D+�׋@�p�+�Լ��h�"�:�L{�,�a��V8�\E�Lo?v D���mtK�<�~.9z�@X��K���gw>g`o���`BP����RR`�L��r���G�*�R��&�G<����?��H���Xq�*TTg�-�oـ�r�t��R�����6�A�$����e��85sW��T�V&*����m�~Є
a��W��(s�)(�p����IP~��( �oG<0`��l��5��,�c.�k%v	����$�j�4`@����G�  �䣓uŁ@��mj�� ��=4;��\;�X���j?�ԪTD�9#��`	^��;��xkf'��9��Ʊ�`B�t�:e?B8r�
�}����)��r����T�p��6_�u���uns\5W��n �lΧGc��~z�~�C�
�E�#o������āS_̢�PP�,��#v�,��Ì����k��I,V���g��5[rt]61���[$�͇�A�؉~p��b���PX��:�:e)�l�̾i���L�5����E�"l��,R�ރ�J���#0.s�ź����(I���g57�X y ����}K�5���d�TpA��ϺeC"��̝�ԕ��������z�v��y*9Ur�Z�9y�
G�t��_�*b�#ŝ��[Vr���:i�LZ��Խ�� Tѿu��� �kl�����*�#	�eH��Ӆ�Kϴ����2$��	�`I�.��o�7�Ld>_�X���t͎m�.���ř��/��Q�2=��'f~��@[�'��蟢��>��)]�KX.�����5)_�����R���Ѡ���X�<n�����,��G;.?�M����΅g6���"��W��5W��v x�<� _�tr^j��>h���:Pi�ܯ����~�¯���v�1�w��^�w��/��$$�޲�>ȩ�c���-DЃ�o�2��"B�yL&⊛����g��+(+��	���|��xf<H8���Ē�$�������@.FU� �S��ՠv	�ef�p;�K�ך�y���6cĖ��E�A�����k����Er�d��^3��]_Ӽ1�&K��wƣ^��Τf#S��Q|�ڻ�^��`j=�4
~�$I�4��	��6Ytvp�L���b��"�e��?-W~����Z�d\Y�FN۩wib�V��Nˡ~�PB����ї��K)����"4A�fK}~����O7��! �Z-gs�����Y����9�C�C�(3��<@T���ؑ�ҵ�f����V�E��}��k��BL(T��u�I���$X'�ܺ��1?q�w�]J�\�]M�#2�m`����Z��1���X`�^�@N5$%� �S3ax���g*�ɆEȠ�@�������I�~p�)�|T���2�C?�������㢣��^���x�Bcܚ�n��΅�3e&��"od$q�3 l2	�Pzw��]�ta�9Nk�"<�>;v}����u����a��ֽ��?�6] �I	u�*$=�ى)���yuO��\� �cw�/7+�6%���������%�}P�U�t/�F�l��L[�$�V�(����D�2�"q��wJt"!�!ǀ���̆8���fD.>:���G�O$�5 rѵT�K����l���w��D9����1�-� �so<v��|\E�S�^,J��]/x��g�K�L��`�Ϡ�jj���vˢD�Y:���)	?�_7r�q
���ah?�r����]���e&53���4�A9�zs+���F�v5t~B��$a���*2�L���=X_oZ�����Jr��4�r��J4:�N9��D߾}��uZ'A�=.L�9?�҉�����[xT�����>�DSbN�+�zϧ<P�\�hO�~�b��@�_�V�э�f)����3����Q��-��	�,��UF�zh݊u�?���6�K"�93��-�I���؀�,�%3��y��4Q��a<E���Ct��ϲKYϚ�1�gb��Zx/ލ�g��;c������Ք����%}� ߿<�����l��(���M���-�H�L"�!^���_�����X[�x�m �/n����"������^��Q8�\SMp4 ���)h����a�D3�Uؒ^�ҩ��)��d�Ҫ�<�B��V���sk��x�{.%{�A�}��Y�pA��b�����&���"�ƨp���N���`ps�m|���˾xu����%/�2b͙�O�~O����:َ���S��oN9[��:��S�G��p�Z�mßs���QXK���m�U���g�@ƲI�[���}ވ�+}.����{9ȑ�1v���[��A]����7�|M�~:����c�I���o�m�4u8�4 c`e:?�4�n�d=�c���/�\�6�jɖ����C!��j����M��OW���=���a�I;%Ѣ%2{���za��ɦt䝼n�h�k���gy�Ѷ�d��i3������6m�[��q�&qS+���{�G�D�$�,�ZS^�rF	K�tV��'��l�@O7�Y��y����+EWɘO.\��f�Y��7�-e��_J�~�96�MΪ�˝�� �v�y� �$�/o��!uP��t]6�lk
I���D���ϐ����M�bc�r�:<�3��`�Y��z����Z��薭��WD~�
DJe,j��j��G�X������	ٽB�����a�+p@S /�U��F�&bZ�*b��M��/�i@��/l��m�M�ү�[Q$H��*����A�*p�~5tn
fY[�h�24�)i�d��ˋ��D�w�d��3��{�a�<3����윬>6���E��CY���M!ݩ�5�<������=. �8�J楾��`)�n)M�|d y��&�^��'�@���&z�h���-w�ypg�c�L0�M�n��`�*
sC�}|�FX�����Q@�5e�F�@ ɸ���l�*��0D���*/�c��x|�%��z�8M�B��26C.�چa��J1�#���Z��t�UJh��)|������4f�i�?l_��>r�'�A+k`� �������Ӹ�y;����2���c�oE6kx0�FmQm%����ȍ��+A��h��p�6�(iҋ����p�k�غf�@�='^�iklp�)�W�}���^�����OC�YL�u������
ɋd��[�\���a�����^�;@�
����ޘ�} �]^�T�&�{� �}U7����Z�T��GD.GT�Cࣻ���
K��%rѱ()dniC]0���x��w��r
@���H��|�E'>����ZQ��69(�>m�S��d*{.C^޵omh���6R*�zV�ݼ65&�G��銙,ؽ����K��du��&߽
p_	��}�R����K�?rQ�>��BS�8,��O6f��FA�"
�oxaiEL��o�i:"Ȏ�pX:0L<�VZج'ع`��+0����E��G�Je�+��t���kh�	<5.�����^�|�������A������އ ����GH��}H)�%��Юc�A��;�Z��PHU,X��at� ߸��*�)q8�	�͆�ۖ��	֩��%�dA� �ۼ:d�'�����C��oI�W�Z��h�*���H<D�7��k&���!��U wj�%���
�����b�g ���o�:6Tnt���:�x��������-��w�p���/3��Mݖ���C
ʔkQD8a�IE�0O˧YUC�-�Y�u�� �:�F2���>MAD��}?0��Jp�J�-7���shG���ڇ��l�x����+Hƅ�E����~t�`w�Q��O�s�Z�)=����7.�? ��D߱�K,6ۅ����$�/�pG}J�ҭ�aX�ʫ-�����OI?��H��<T؜�(�_*d0l	�L�0��n��5o&���x�92����ܥ,J�4v�5��5�y���+W~\�ir �TK�>`��=Lq(�*��H/��'=(��ŨV�>J!���&���}=*�R�'�n��������z&���xQ����Z�^��R�FNё�}Q��E�pZ'��#��Ĵ@�tf��mr5�J��O����[��zĿ&�5�i�������Nd	2o��K/��v�v�P�#�mt>2���H�KR�*����_I?< ���z���	����x��x3��"9X��>��qY;X6l���2��Q,�a��>c媋�c�25v��n0cI�<�K�t�c�I$��w�ř��������_�
�LS�8��\�xd��1}�K������D�E��"&_�4$�[�Y�z�<��իn�,:��`���n��E�((:\Y�L(y.=�bk\���ȵֿl W{�V^��@�'����:ǒ"f���bW�����'���zÂ��>70�L�R���Pa���N��@T�&(��Н}2��\��������3��r�SO�]��~�yC�(�h+�+u����G7f(?���+�6{�
7�GyH��Xy�K����(6j�ͽ����B���ƭ�R|�������3}�����U�43"��Qہgsij�T�h6^�Y/������f:FN�^3	Pw,FΤ]B��(��	)p�ڨ3�Uu��,$˶�T(��^�Z��_�f�@\��oK��l2.Bڋ��KX���и���}UDc)A7G�����2�Q�i��b��|`��_�{z���v�"��ϛv�m���$?���^�3�Vo�>4C������ ތ/[.��+j���x6��+|�J~����T.��
��[1T)�C>���}�J����w�inw7�f����@i�>|��p�F�*��6(1�cz3�T��J�ل���U��(��3�1���]�j��o]pc��E8~�gs�A�x8 a�h��աD�e���	�,Lb���ԪpL*v�-x����J|���g;��~�(�t* �}`6��S�������D1*�{".��Ǜ8dp�c@�5��;��������ֹI�a�8 �&��x���h)颿^@��h7i��$١�: �e��*-�Iӯ@�?C.���(�����ҩ��ObLrh�n�~���_���\eOmh[t3j�#Q�mjkS�(�e������8��Ng���K,дo9�ď�_Cw��?K��j�1�-X��8E�q��:e��\���m٬}�������,�xz���̌^9����v+T3�%���Vp�����c�!���(��C̆���K���I>I��x	�[Z��n}�$A�σ77Jxް��b9�#z�=�I��m��7u��s:�h�a�K����k��h`[����ܝ�Qo�$Rv/�f�#2�1U�X<r���$٬m1Xp��G�A�4KX77Yh�Y5��O���A�,�w��ך}5���bF��F&�L��jSl�z��}��D����/Bf�8�ts�
�(��p�	]��`�
���)��N�"-H/�"So�X"�%�]�Aۣ�4��z�Ecg�I�}�A&1�M��/+M�fԀ�M.D�6��_g��3;`A�w]�j$͟vAfT7�1� �p��u�$�ׁ�8?�t�ɂ�+�w�������.1#n�4;��,�x�� 6j��Q4�����O��%�/f(����?�#�ZU~|��X�����/����VY�Hjj��gK�`���8@�D�f�j�۔[J�����˄�9:S���� yz�����O\G�[��.1w�/RM�ԍM��[3n^�$ߎJ���|ZrO�*	���	���djD���h ?��m%��fJ^�r�>�]��F��	OwcS�eo������<���\��E�3�͟CrE�o[P���F�I�x(���p���-4$�)����;�P�M��f�䑝*$]eWb�G.,�e�^�Ah��V�Z�V��r�h��_�r>P�i�E���#o9$��bp����m���S�A#��&��X�o��6�Γ�=�6�OWӽ���! �L�_��Y(�^ q��ኰ�9ӌ��DY(�V
�̶��^nA��A:�����;/u�=@4.�j`e��<t3���l�Ǘ"���MJZu��]��Z�SA�ye&�LV{INg����.�rj<�}�� K.
:%v7a�A5u`�$�:{T�V��$n������iل���~��n&���W��e-��58L�c�l���b_��̓2�9��ѳ��rK�r8��$��艠��w�$˸[�n9(j���E[e��+�ι���V�Ļ�n ��Tz��5�s�F0]�EXh4���>���w$n!&��?A�0B٤ý��et+��O�X"�(�ԉ%���F`� e[���R�����~+vS�]��,υ�'��kNx�3���=�u���VJ{��Z����������?��(�/&r���''sW�?�Qx3�e��N�^5��^k�4�e�k;�Rӭ]3l��R�Z��<$�2��ָ�Z���3L�<�;���5�h�?/m��/	��b�nm-�Jx]��x�:u�vF��͞�r��	w���~�ҟ�Q^@i��`���~��JV5�+^q�ge"˨��"�]%�%�y�^�q���n����Vu@�����9gV����*������x��h���Xh����͊FgV��;��B �>R�ԭl��
㋡c;�E����N@�E2b�F;���<q.̈́[SE��/O��0���o|K;��� T0�����P������ѹ��4�����ֲ� {$`u���r�7��Yf�=� @�/f˱Kz��9��n�{qsZ��^ЮuD�.�Y�zRn���R��<9G��V��v���� %"MI�LK8�I�`��o��BK9���ѿ���TY�}$?�0 1j�v��`R���i�1y<����Cw,��%զi�]���H��A�7�^�_�8��:�\���S��n��܆��9����?yR��׻X��!A�}pm�� db��p��ts(�-RɈ*�z����������
@�"�H+�N��A�����46���Q�L��!.�`�����d�7�"�n�(V���g'��������[ȱ��
>|%�S/�~cP����t�_��!�k�H~���1��;"s�<f�dKa�4⿩��?]J?��` 0��@��ӻ��]�N��L3d���{@Zu�i�?�W�L/�*S!
�?3�%M�lJ���_t���+鳷VL�
�*��ss�Hz������9
�I8�a��< ��j���;�����]1
�O�8��^q͈	}t2�*%�W �J�{{T�L��,?��`�����4�}g��HXEx3"�6G/3���r���Eã/4Q~`�c��	$
,7���,@3�H��s��y��c�6������Uoi塀�,����
S��-"��v�oa�	f�r���n6[��� 8N�݄���uы��lC�ik���C��#�&�VP�h��<�0�(��7������Zg̺c>�T���bz��=�u�w�?�?U���W0�?���༢��1_&��)(x1V��C�E�I�=���DHUlӚ��@ac�v��������KҖ*AB�X�s`�ͮ�
?M	-'b�Gp]d�(6Ș�%�\�γG�Ygs���O�@t;�ႜ�{n`�q9w7�unbf)���mHX���/���W׿@]�&���,�����Ʌ�#%�-�$�~-�{$�7u��i�@���1�����Ǣ?~�j�����e&�O@�)|K�ݽ�`�pŁC��q�Jfe���I��y�������)�6�ď.]�O�P$6wHu�=o��C�g_�^��D����<o9p84'�P�Rwe��jMB�Ʋ�a���l$F�#~4�����"b�Ö4T� ak��8,@Os���zٓ���(��L^�GM����Vܡ~�@c;��"�jp��z�]����n�Ĉ�IrH2�/�����#�i�5����𙔽�2Ub���E4��j�J�����c,����
&�5"E�ٛ�g_cM��P��_׭]�	�^IQ����x�����<(	x&���π	��`z���ME��?�j���G;e��_���ӱ<��;DwUz�n U��2�G��4��g�x��0�$I|˰,�t���g8<������}9`�A��x����هZm�.�3g�m/�* .5j<��;3Q��D`���*ݡǇ ��2�(��_�VR�������a��^tF~���~��:�αT��4P�wC?Q�[kD�]y�x!m f�+��HД�*�83)�s���9��O,յ����1<-71�Vo�]�`���
�s�	*
Cƅz�L��
א�V��U����^L�)��00�R�\zƂ�����BѾU8M����m�>$��biΣ�������ߞ�s�+�< �P�
.ϡ�T��sC8m6-�0ҥu�Nw�\_���.���Nk6�ܧ�q���рO,�B�:�ݒ
q^�W����AΌWĎ�����oO�a�x<����pO�챼�~|���s�V`Ia��Z��{�_��Ye���0ϵJ�����$9!���Lo�[�Y(��Ú�S^��y��Y?�9J�.�,9��G�&��Z�B_b?�;��L��A�]B{ݞ��8w/:��$���t�K�2Y}GNX����,��H?�O�X�P;��h%���@�����[�"�X�E�+#PhS���'�6�Wf�Q���s��mS�����Bl���/���Gl!�q�����>-A�s��� �g_JZΩ]�/5/�0@^�B,�Xq��.'w��:�ctM�w-���#���Զ��c<jrl�.S���TZ��qPl~���J�tT|���^�BD:a��CkB3����&�97�$�mT�Z�V�U��������3��8o�uT�"�s�������>�{��U�.�����[^��ßw���� '�POG� v�-b$�҆��i\X:.�	� ���)��=O�Л��T�W�+�$��l�s�aO��I��rX����-�V���Mxw"�	 +`;G�i�z�`;ϼ���,M�
$�^}���B	T>��[ն��̵�=�(e
N[4i�0|���ً���O��� �b�9��A�$j��^Y�>0��
�ԀҔ��'���/�K�	���y�c�����B��d�$���.Դ�T売dX�a֒BH�@�����{��D����s�_d��_"� x*X�{<"2�~�R8�P�3�=X�"��LԬ�~���~�
����c����.�},ap��[�����!3���Zt�,�PJ�P�W�*��K�c֘���=�U��x��xT4��nY�,�/p�G��5,5���<�6��Kx�
�{�S�(��-Ya�u�x�~��I-A��؅��U�k��V0�s���7�4��������:h��Tkj��������	�]�=�{��X��j/8�^MD�x��H5��gRj��;U�E���qjc�d�e;:��:V�@��ؐ�������hlcnK0ݲ�ٲ!ޤ�:��B̽���R�A�y �^=l'�t��9e)�IC?�'���� ��_9MF�W��W�h7�5�\�DYg�H D����Nkf��خ5{����	V�uO��N�����<%������x�I_�r?��|y�t�26)��G#�C����	���n��P�X���F��͙���
;Ν:�,^�I���4Pø¬��'J�d��h��u���*��g�%nт�_�i�B�C�Mʌ��7�I�h�KWsɰ����1�zF-�k�}$�p�A8��ʥId1�[��0�9l�M�J�C�D&��ie�����/hͰ���.=+~k� y��	�k���j=i�p� V� �:���"��B+��^�W��,�όu�(7j"�(8���ϡ�3$���ln�P�!Wʊ�;p0.��&�!���(8`!G��-D�-��=5���62C��B�w�*
��PV�wnï���5B�Qȕ����Q0A�bxB��X�)�}L�t>�e>���@ʴ3q��/�r�vҥ�^"�ϴ���a���v8�\����Y6
;o�-��r�����fW��Uv��3�f���x�V���lA�=��Ed�	�#Kg@�Qc��Y�K18�
��Úʬ�ځ� ��PX�u��#xVj:g��|�<�i�Y����)���U|W�'�1ݥ�4�Fx�����a̒�+���c��0?�7?VD"I�6:�{�ܿ�1�B#��m{G4�,L�Ɯj��������w�W��ԓS���Y���b[��~)��R}�fTv���+�[W��k<��	���(	#��j1T N���HkL^��I ZK���\i�2��~^�@E��7��dٺ����� �"ęe��~�5�iv�o~���,
��I+�XY���q�����jhb��EM#��C%T���82�uP5]r�vQ�%]:�ޑ�D!����#��S@��Qx8�:�N°�����V�}����n4�}��	�����Ҏ��k�Ɗ�+y���.ɚ L�~�P�9��z5B��\|C(�s��}��f�?ϐ��|z
sKi/B�a��~Y:�k��n�#3NsR'8�U׃Ą�"wrgSw�%����#��/>�H��^�g%X�=�ݧ(8T�R@�9����5��J��V:!�&Ei�۳�IQ�"����Q>K�)�}��"�ݨ"^E�2>-�x��'�;�	 FδCش��5�-r%%Zt�ȬJ�,��>�>ژ~0Q�˴0#4E�W��ڨ��d�3�ky�Q�(nTH�%�� L�z)n��C��L�,��D}<L#wŤ�����e,⢜_U9:�Iģu���!�dz�x��)�d���y1��U��o{<`	�'�OM
����*�0#'�k�,p�5�Q<��i�m)c�>�D�)i�6X�en�6���\�~4&�s$�Q�6����mz1u�n8W;be� t��{������l��C薿׆�" �b�8O�6! ��㖎h�#�����y�3��EVl��l�aE�������J�d=0������A˞�uE*#��s��əC�Σ=��2���Y����A��.�Α�.w�w'�G䅬�����������%F���IM�ȴ���ş�lQD�xqZ̨�yIS�x�6��q e�;��	9�w)�[q���aY�<aR:N�a7D��%>  h聎GNV�2����w��<{��gۈ-i�ŷ�����EC�NCD�cT=���V����2=c�lYQ�B4�a��;T��Z_�͖�c#�����.d<`�K���+,�뿁��_Vͷͭ/9�z��\��w@���j���v:�����Eo������6���hg7r�Lα���
����%7"1 W��Z�����
��c�s��t"�*Ү, �EY���?�vk�m�;�!MK��\
�&u��.��L���c���Lj[��&T���+[6!:dMYಳB
z&���x��J-�QʘU��q�u�9e�f���jtiX)��?	��g�ԁ�2w
z�5Ԑ���Y��E�xhښ����?������Dq[�wf�A�q�]�:k|�Wϵ�+x�Hs��!ͼC�(�Y|��琓*�=(��A��M߳a���x�z�ŕ8� �l�_N�4�����6.>ZҲ�t*Z��~#-�����e(�_��.*����gfX�	0���/�79�"����z�{-�sB��b��<r�>љ����ό7�l)/�#��=�,�@�6����5P&�����^�]��nk��:�s��Q	��,s ����ê���|�N�x�\����/v/w����>�ы7��:�9С�K7�o�\L�3[�Q��TP�2O�J�P$�Ԉ��!÷�Stҝ�|�I�� �y�L,)A����.8��|�Pfg�#4�8���&��JJS=�8���#!�%�U�%��ܚW��w)�m����p�څ�3ݸF=�C(_�p��ץ����2V�I���� �"��L3z�A�tY�a�~�c�J"u߆Xfg/�Ж<�
hY1b���M��'�}^�:����r�ؠ���2u��F��$��n�hmƺ��SCRN�j\���+�:�e@C?f>�ۉ:�V3�ǽ��6�d��?�h}h��>V�B��� �����B*U�5n��s�8s#�*t��{*Uȗi݁w��`6mfx�Dn�'�5�l���vR���a�տEv�v,�Ra(Y�Q	I�T�D8�9D:��oZ�)����N�y�
ᘊ!�O�x
�UpہU�{h� �كN\�C����#.��k<Y%�._�펢��}��vM�}��l��+a��OR�f�H�y����kĪ/ :���|߬�!��W�:ѯ��|�2U���f�z���خ<�t1f&�7��Й��.� _�Z���C*z|�8ޅ0˧a���R����LU��O�7������p���1��m������
}�����P��d
���ka׵_T>���q��Ѣ����L-+
f��]� ]�dod�߈��l
%!§/��_c��b�tOlTѵEт��-4 �0H���-J�5U�P��w�|P�o��1&���)3��ZI�du(��V��D�×��3��=������@m��ޙr�T���_k+��k���L�kC��|�z�o�8|�gݫ5�b%^ꮩдH�%P�ϥ�R���{x����|*9s��5R���C�#�b7r\w5'�>+��=P;�eS8���cò����D*l;!��ɺz/H�X�xxݸ�El;zW
��A�(T��̗W �����]�4)�m_��Q����T�U��}���}d^g���&fћ��I���!B��+z� +�~��D@%��/g���W����7�wBCT�.�(�H���؛�ȫ��`X�v���6����u�;	tFKq��P���mߎ��>o��M�� Q�\�c)���HT��Tl�����n�"et�e��!��c��G��4I_�XW���M�7�7�϶2"�������[֊ϰ ��ѐ0�ޕ���3���=�(�Qt�c�!&�6��f~UY5�F22џ��p��|ws��
�?K�s�$K���~�{�op��܉�&K�&j�^)�u�m��˸kic�ac��:D5.s�9V�|�޺f�z�r��H@�(=������� �
��E��,C�+�7����Rcr�;��i�ݣziC�`�
r�ݳ�h�1������sU�LU@�_A�;��*z3yd0"ͨ񗈺��ډ����������{��9���k:�#kd'd�҆��n���2lG���j�j����i�-��v�Ё�qI�����v�`M����١��2�?��v�Y�e�1������֙T~���/T/������"�z|���ۥgߒ"�I���wiо�=����6\3�����!�k�Ӗb�]�$Z��rB�VS�ns������M"7ѿ�T���_���H�Du��c=I����f��}�ez�8GМ!g�tH=����N��|D�����t ���@���k0E��WW�)@K��Eoes.��{�_��Z����'/i���W�����r��1�:�
]���!�Oz|5�.����O�9]�k �j��XZ2d��D9A��z�sLk7T��c��0�a�7�"V�i$����X#� �ՍH�eW������/�gыN4�clj���U&K�0��B��-^
Gu�#�X���t��<x���pc臛ҿ\�6`b���G��ZĄx���[%'��#����[L)Jز��1��`�IӧP_��@BzS�Ht{��R�%�8�[�T�q�2�R%07n����c�S[���%�h�eq[�?@浈�~������?,�r	����m����b6г�~�8t}�פ&��3&��vb�(�(a-��p{=|��Z*pG��a��g�s��\�U>�����#�-oI���P��R��H'����Hֶ	�?WX�w��w��Dh'��;X\�̯cf����q���TF�z���� g�1eʹ������R�;V.T``1,$ns'=9�� uQ��F�E��!��Iq�.���Jؗ�7�Ct�, d;զ�@֝����l�C��y.1��%�����5��|�ꃏ�+����Өک�d�k��������+��SHǌ#�G8Zf�)mA�3����ٹ��mv�hӰl��J�Ӓ�)C^|��3{)IgZ��Y2�5�[�ށ+a�}���{��d�?��3���a4ҝ��x�l�x�9�P�p���g[�^jƲ��\+u�W�.\8��k�"m֨ZF�3�W<R�u�㢵��r+zETT-���Jڅ������b4Pl��O�/tp�����������,�<"u[�f�@�U�8~��I"�;�����s�/�e�U��}�+�KㅴY��~�.ߎ��#l�U�]�$1�.�6���[��
Vp�V�W���{ �0�Tj_����ɍӖL~���5
y�oZn((�%c`n������lJ����k�ĪG��*�`!ڮ���i;bk�Y���3���t	�>� %����%�qIs�x��E�L<p��� �����NƆ���.��9��D�eįØ�D��όI��>�Q��@�=�:H��-��
���}:CF�$��ܧ�Hn���?��GSa9]������aX��P���Q�-����<竭N dvMg
��~E̗c�2p�Y�u?�XoR�P��P���k�e��VY��Vp�s)��Uh�Oo�Y�\���� *\;���q�ټ��(E�&,3�0u+|}�����L
=�\�Ma�)e^�����·<��ݲ�ή�w�q�c�gC��Cޅ�g:�w�?�U�O�'���x����[����z�!:�f�`�nŇx� ID�`�|;���b�و���D�G�u	����6,�,<����9�"ŀ|��+u�2�#*�*-�����R�Ř���F�gO��F{�Iw�����񖐸8�����D�t�fW�I�&f:V6s7���_�Jb��tpw�
����Z�'��������rN�K���}�z�y޻�1]U"�$��6�d��:(R���+3;�Q�uԿ&w3����1Z?�M��7�I�*�eU��>ّ�Fh����9�x�>K��Ǻz���֪�&�<�X(L黽f��w)|j�֩�~	�e��e�*��Ċ�g��I�\v�{�8&f�VE�^�^��ڈ���;�_��.��%x��$!�í�'e��=w`�/T1�bu`�h �wj�l�RYj?�^�Ȗ��4I�1<Jӣӱ�X�\�
6�vH�K9zC17�͸1>�A�wF��3@���;e��[{U �ޗ�	������p�Je������>��S���g��/�顆�[͍e��X�~s��x�݂�Ϭ�/,rHt�8'pﻖϠ����X�r,_�����l��Tg���BX�O��L�z��0'�1�i�ˮ�@.<����MH�^�}�fOm�H	�����7w������so��R���pI���z�j���Jn�bft��,��l%����Km%eG��,L����UU��$�Qk�D,�m��W�t1�Sgċ0��!�#*VRp����6j4�y�o��2�]�G0��=�D`����6f���	k.FC������j�
��__V���&^� dI��}C�@0:��l�v?���>8
�9��:�%_�r[�۵u�t5=b_����ѐ�sۄ-׊և��S��;��1*��)�$�!+B�gXzLc�yI�N�]A<�EF�y~��/j��V���;k��g��=Cu�Ùs�����W�h]笅2:� ��c�DK�5�{AX[b'I�i�t��f�Ȫ'X�sd���#x��8���y�^�w��EQ�"fv���D]��P)��`�N�mH�E�K�Ϭ�=�L�0"�ɀ�9��ޖ�����[D����"�����ud�%OzV��yn�d�u�_��|�X,�==���d�8y�h���lT���
ѢHѲ+`���M=�MS\���A�����ƋB�N��W򦋐Qb�M�s1�|��Ӧ����j%���
���A�CF���Ћ�A�U`7�(��N�M�)��x\�;��"�XW�~�����ur���K�{�ue�4�i����0P`]̜��uz�ۑ�Ƚ��V|(-'B���u���m�k�l���[Y���Jm������hxp%���8��Eˬ@̫d,�^<j� �j�ȏ�#d
{�CcY�z�L���˞��żW�J��]_��$K�`Yc�G��%�R0���#`�¹{f���d0,O>7LX��SV�JN�����h�^�L��hlQj�_"yq0	��{
��W�,z;p���{�m�g��s��3�E�,
fG��[�1ǀ�fr;�����'����R$�}"9~�F�Dβi���U?���Ҷx}#����BY��^g�����ޛjFl���xƏr��h��G�#C`A^����.9��6����4����{ӹr��e�/��
�2��b�OY��{�7f�n��K�8��y,^Q�3ֲ�i솳�D9�n���z���nl)�����*/pbĎ,����Oۺo0
�I�U:8~��.�媭B�q$�۫�(�8�?I��������|��s��	�R|m!��!2�X��M��,�͟�e�UC��ǇZ���N.��V�^`^��"|�3��4j����И��GoS�	�]�F%F 22w(�ΠuVt���3��va�2��.��ˌ��(U�7����������
X��=A[iBv5&/�~#���j���%�	�|�b���JԽ)��ó<��26�)N;�UO�$�?{b(T:
����Z
3=��0�{��E��㈤V?Ck������/�r
��|����7�bT�ձc�!r�seI 5V���Kt�9��$����r��=���RY[��Z���tJ*e]`y�5l͗Ү܋ۦ|;�u�k��;��jn[��+�+�v�$��#@R�m�[��,��dE���G�Y���.|���[*�x��w�~�Z~�1��p�69��J��#0V�nƄ���c ��!'+>}�^�����L��� sn����cP�W�;XU�\�~�=�.5��5��g�e~��UE����`dB�N�.�e�P���bs����Z�
�_�p}�!�3"�]�?]'�dnBC�4EH+�n8�%�PD����q�]�r��ٞ��i�Qԛ܌����m����V��U�MR�"h�C��j;)�Wp9|��L�̖(yx��v_�b�CM~�����m���'ن���.�n(Ȋ����]`�y��/�Q�P�q�F-��XD��/O�{�N#K��g�5�=H�	���D�&�d�p	����!F�^�l6z���ͣ�P�L�4���Ak&W�����^��j�,�D�UE�&Fg�D.�0��F�v�=�+�1X~�$�ؗ��X�T�+25\K�a�Ϛ�H�,&�E�ao/�O�����p���#y��/�o�����<=��V�B;l#`��x��5�������{O��A?����i�4`�*
�Ҽ(���g�I�`�]�>� �F�q�g<ǝzQ����D��7�p�� �}�� 3�d[x���v��DT�O��b��9�t>Ӹ�H�RԜ��+����P�ua�L�r��8�/⥪[i'l{>�ט�?y�����$v#i������#���]@#��r�R3�(�`�&;��d�nȾ[�P/iٻ��v�,v���R�Ѕaw���d~C�A\L�Oxk�2w��Gfa�;;LZ�_���ץy�F�e^��cؒ ���`[��c�!f�/�%�tJ�(�i䝾;��.�m�i;:�E,�JFɰ"@C�@٥n�ъa�a��Ĵ�����(�ڒ�����=�F �b�o�e����׼��Et�d<&���,lr�X$I�K��B��������%�(�����~�:5��)���8dDB:w�K��U��ŭ���g0<�!��|d߿ZE*�9���7��L̄�1���_Ç�Z���1s���v`�w��0A%�T�Cy,�|�B*'��\�G/���<���"*�����Ս����c�Mnk{�:�D�����=h�u�LVp��p�x�qpӵ�R��	٢)�۲&����1.PB�~'Ю톿���n[���p�U��z���gvK'1�����FHѸ
nf�B�Eeج��,�X�{�h�?�X�&���>*U�)g���H��K[����%�rI0M~�:i�%�S�O�H&�/����:\�kn�E�ꔂ���M��i_$i�"s��R���!� ��4���[�M9��^Ǡ7�(:�XO	9S�b�]�~��VqD���ҾS��<F;������p��Ŀ����Z�KNe�Pz@ݕ��R������ Hʪ�L�{*��{���/��'$
��m��Rp�P	�ŧX
�y�Ƌ��8�ds�SKeyT��ɻs�״{��z��{~��x��a�9���*��kbR&=������x�9
�_t�.��N�k[�.�d�ʟ�?��~�\������)>��0����`Y�3��w�Y�����a5pov�y�'cD|��a��W�zrc$*�\@�?j��Ki���b��8Ͱx�ar� M�`�G�/�7��\�<�l�%�6a�Xl~?�4�9��`��20���;�߳�q�M{��(q+^{�Kok�^����� Z��������9���xΊ��0���d����Cƿ+��a� ���&�p�.�f��բS��0��L�k;q�lZ�8*�aɻ��}�G�.�C
���ӧI[�5��Q�Y�/�\���6]z��Mby-���,ʢ	1):��)�{Q��4����ꇇaXQt)&�3ݙ����b���D$�=h���7�t/��v����I��Gk�ց3 +�t�C?H�a�U}s�T�z����i��N>��\.��w��Z�������ձ��k���ɳ3��B$|�i��S���o菏J�t����[s������������6$���{��س�Zs`�R��@�$�;_���stGm�ć�n��O��L���Iwcr��G��4̽��!��y�ꓼFr9N�����ߴ�t�'G�H�a�{z�wh�G��yCu�ׅ��e������"�Q\4��V�(O���[����(4��P��T�n�qx�t�g�i,m×�sS�gא��o�i3o��u��V�|Y׃������fu���������+�3: �>�JD�^�WB 6П�aϴ�ud	[ ��u�
-nV�}A=ÛO���D�o�o8�X�L=j$��
3�Ы��|�xj�`��|�f&6Q�����[r��7i��J�xx3�FCQ�Y�?3Q4Y	G#����m^���ǌ��vИ��"�,��i^�)e%�k��Z�/C����8Y���-�%����s��Ҟ�/�D���5�=�{���AĩN�L��/��jȳ(=յԂS��)sU1p��a��r4��(�@��H�q^��mBei��4�V7��a� �nT��`��C��98U��+E�>��tb��{j7ȥ�c oti���Q=����V)^Yoܦ�����\��L5���<䅵���]�z�C�( �3h ���.i�3N��=	�MK�Q�iLP7�K��H�_}䴐tͿ�&�R��3�+�D���On+�*��k���OӞ{�_��"Q����xH3�SUC��F$��'oz�f��O�B���;X�������G>�Œ���7��/�i�q��q.�a�C�8��
Sk9-���~��U��b��V2dJ�<<X5��H`$]����C=?�������P@�Ƨ���!k�Y��N6�U_M�u��W�=�RC]/le���]��Wk��Jg����%&�[�|��ct��!�P��M�dsj�D�Q�[]%��Z���I�:��Σ�轿��X5�+�a$�4Ѽ�C�]��WhӮ��b�E��>$C���Źp��3>R*�� ��hUX���ٽJr��|��\����p�_�������񆂾��Ұ˫���\-�`��-����{&tyX|�G����#��ϫ�o��_��P�)��Z:�~BR��Q����Ak�m_'�e4���L����f�W5�Q>���	=%Oh����/V�׍�=��h�'�ySv,!��HO�r��.X�������u��}
�K��E��D)��N	xD���X��M�fM�7����Ŋ�M��i#s酁/�$e��=f�e�ZQq��u�u�;�OQ�]�<�.�$�
:���|M�d�<�����՟Y�p�x�7�e�n��-�������H�|�%E�b����~]�Q6�˳��$��}����)�C� ��VQ�4�e�%���^e��u��F0��%ʽV�F\��0[��f�-ᨌ��Y�Ki������`��x�~�6Gg{�����ub�@�;�U�Gy ���)Xm���J-Ժ�]>��.(<P��'��	|t��lB�2��������p�i
o�*"ULF��!��B���oB[s�Z<m��ɪ���܃qUC3#��gPbM�S�9���-���Ps��h���`��Z����d����$" r�l~"���O
��)W�r��d[���'���I�_D}�Vb5p��N8b_���mL!���)訖�YN��֔�|�F��G0�C���P��l5��l�ƟmD�ս4v��#����p���P�Baf�{�n���{=Y<���惜�U�G�a���lI�x?���p�n��~����{��`�Z�#yb/tA2z��4?�R��&��eʏ�{��+��%��3�4��W(:�%��^� 0���
��0rYIF׾\g���v��1��~��ȂfІ�Xϫ������p+آ�!l�	�f�A9��^}��9jmUT� ���ϒ���h�xw��CS�
̪m�ŷ����#6��ǥ�F�γ���~N^e�Q���� �!C�x�x�z��=�o,�W��G�	��9�c=��T��J�^bw:%����/J�%�g�:�X])�Hey���Gl�'�Kt3+T[�*����t�:��K"*���m|v�b�[���Z|�EōkqR-���:�[�pB����\��>���l$N6���7`�c��,�%KҸ9րbb�c&���ڲ��>o�h�͐��U���J$�~��H��,#��,FR�f%�m����m7��B��Э�h;��0�;[d����7�S�s�Q/mB�����}4T��7j�B>��7�+������Q� ��������t��
^�Ԡ�k{�>D��Z��~����9k�]3��u�y�+-�GU�h��6�7�0��bI�ꕛ}Z���o��o���hh2֛���x�4.~�D?�KDk��xH6��G~�K�$w�K�O6��(Ph�mdj��ڰ(���>���+�l$Ȟ8EtnD���$��x��N����qJ0���ƹ-`љ3�?y�5F�x=$�d�n������ 0�(�K�c�T귣�5����:�q"���k��dpg���`|�Cp��ϧ9eB��r�"�#���1
upr�<_;j���L�~`é! f:4*vM}�L�����>��c���bd+�h���j�I��m��e�� 3hzFWT��/30(fz�K�?����	4�W�/t�6LN�g%Wuz!�-s�ġ��b�в+i���AQ
���F�H�R3W\����;��S�M������[��~W	��s�%�����>��Z-�=��'T�T/H�[��3�hשIl�ȯ!	$�1�����ITq";�9�ʀmn=�Z�d�VvY {�'���C����,�����\�������tU^JI���:+(R��D�dd䔻s�+�ڼ�G'4m���ƻl��*禸x���|�F�����Ɍ��W!ҩ���&��������M��6���p�8����Vd��G��q�0�B{/�o�22���� J.�d�M�f�L<]*fܭ�K8�Q���Ȁ��Ĉ�����v�d�n�z��CXz��Ȗu�9nTOƭhjj}�R����L��_�����1�p�UC�_��b�H�J�ژ���jƯW�1�@�a��۲�Գ�TvC����>�2��h^����L��A��&}0�8&.�ǥ2��L��\y~zF����MJ�t�G=��&�3k-�A��m(/{�Rc0��w��<������_�1\t։��Tm��`$ґ۶$/�*�l�����`����'�d��%FP3�ǂtd���դ��s$̞��!^Äo;$�����6Ѩ0�T*G��
_�eY㊕��Y����_����=uFx�����Ij6���h��ڗ�:<��SAfwQO��\��U/��t���d�Z��v�d��@E,��I� �а+���l6�U��n��Q�X�u��/TĬ�_����j7��K	S({������&/�Z��k
���a�k��e��+f���
� �v�s��HWP ||֙^�SKn���1�]����� ���M�A"�	b��_Cݠ(���~>K0J�5�~A�KN��)45�Y�*����#;�z�R�h��m߽|-��=���^^�[��<[��Qc�s�w?�C�+Y!e)���e�����a�cN�#�>G��[�=�@�{K����DE��W�ݲ'���Qm,�۞�"P\�$�����Й`�S'�G��^mC�~L���	����|�B+0�[�ә ��zk�0�vx�#J��i�c���Ί��#2��9׊c�oVb�9��2��ܻO�!����/��xX�8\��N���|�(�U*&٭�!��e��і/o�)!"G�E���3�dPrvE�Y���9gq_=Qc/�pv��Q%y���id�՗HƍG.��:[硒-�ג�G幜���p>u0
�i[�.QK��_�=�R�eV~-�Z]3�_��fo��G_��&�Hr?.�2%5a����k[�E�_u�	h Zï�^k�FEQډS[��5��� 	��3�!�k-#]U��4��1�d�A9gTlʨ�n,��+?��(�9�w�jE��x.�"wS��o9�~$9~�C#
��A�S��mQ���V�hI�����m;}R�a?�d�����E����µ�!��
��}������02�B[D���o,�e��W�&����P-��A���D_'h���H�Y>"��f74�JD��6$+�� ��t�3P�Ʋ�z�CTL�6vek^*�ܰ���)�UJ�=��d���z%S�E��o��N�c FAYr�/YE�i������H�BbpPM���`H	�Q�.��7�`��"��EA��c�|�"��~fz��dNWxY��#�`d`�vp��(��DӰ�*��ĴBI�b��}F���[%H��b�u��̓������ ��~�1�)eNv<��R����r��fJ��}yB��iߞ��Ty1O���+I=|$Ս;��؁�eŶ���SrE��Y��q<�n��)���%TI���V���w�@e�=A;ˢ�k�~��|�8�|7XӕJ���z��[�/96v�(���&3�ӟs���"l�W�lG�h��ю0CBN�:�M�h ��,_�"�jѤ*���MbMNɒig �Œ��It��=����Lm��i�B�5��{\�L��|S�2�l�hI��;0���_@����5�x�5�_�.�V>t�Α��e�	���Q�R�?���a��S}?�t����ae�⾠��!�t4�}~���5/;Kr?�I��3���*�mу���X�}����H�a�S� b<�v��B�Ʃ�(p5i`�PP����>0;�#+�iv�]���$@���>k��0aKZ5�׌�D���^�.� �Z䬑3iZ	vѵ��G����T@9��h�pJ��x���t��	G�mv�Z���],"Ga�ڱ��J��2�.�\
Y���*�q~�x�p_�lӊ2r7�B�2{|��{�י�b��1	y>�8W�����"��
_��zQ;FKF�����Ǉ�I���Nk,��T�$_���=(s��{o�/o� B�X�>��܆��v�t<��Ř�0��1!LU����e�������77���r�@�(|�cU1=<R8/Zs'7�Izf�b�Hhr��3e����$/^.tGT����s�K&����q������E�BЬ�/K��9�1�M'��i�vw������К�;�V ;�X���KLdԕ���<��ی�:��0>x���z�!�	�U��%DE^� #���_�عp��rZة-)��)=�R�-��Aԇ��9���P/�+����F/�*��Y�����h�l�Tf�8)Z���]|`Uk�d7�(`��T��e��p�?SM
�BZV`��Q�E
�M���]I�g����.|{%}2 �G�w��F���<a�1?"/.�&�}Y���$6��k����*��
?��K�����([ �-�y�@�7�@�B�aM`�o��^~\S]t`�Z8�\5��]d�9���5����	ڽ�K؊�-E�!��ʤ�V���=�h�օp�٢uT��.�7�R�ϻ&��"��/)�������z������d��[�[�a� �߽&v�^��}��$;���v7���hX���
N��ܹІ��y���y�><�Y�qx8Ų��Т�"�1O-�Zh�b�"E�k[��fզ˘Ğ��˲�2�~��/w�e�CM&x���mf,^@�-�YD��4�k�v�r���/W«�DV`�bE�q��<�e�d`�׀1��h��r���+Qv^�nf����5�By�65;IW\����j��9�,B�s����ZڞE���_~g�	���eZ3��x}v�W�܏��ZK(Tr���l����`"�����o�����vmJR�������ke����G��EW��ؑ�g
ntطf76L����V�yQ}�/،xJ��D�D�����.C�\�S㑍����Ů�]i.��p�&�����ZTY�� h�}�l�D���A$��(��ӎ>�^`�&D�t�%���k��k0y��E��Y���I�/dǤә�QfvI�����[�x�6�T27'y4qE�L�=�����q&4�,:����(�#>N,��Z��`��t\�!�sb�',��o����<Q���U�b���p'�S��v������qi5m��5��N
��d0o��L���3=�t0P���;����G,J`��ք����J�����R�Z�T�`lO )GWK�� �z@���R�}O5�K��]�W����K2��lu��{aю�����G� ������s��/��L��[��2�{�X�@A���O��N�|4k�	qܕ�Gd�y���4���i̵��8�Ζ$��XW�	����l�g���˜8����5w��Q1�0#��B�֣T��zi��^��j�'�'��T��pŨb|Q-g���AD��l}2�v@�Q�a��G�$A8ߓ�$���e�E�4��~�0�N��k�X��Nx�.��J6\M�e�a����OC¤TGk.ن�����J	ثjQĚ��Oa�,�s
03�35Zgd ������-�H�0����o���,/��~ٍ������Š�q;�X�0��@O���?c�W�H���V�+C	����5ˊU�4G� 1!�4Y��Y���Q�����.��?|�Eϭ`"�g�2'ϖW%T&�Tq���`_��3�����oVz�o3��Ԓ(�L|��J���ʩ�:��9�.��鼰[����X�AphY,e��y�F�ݓ��(�&]���=Ƣ'��,���:S�ё��\�7Qr��~)$P�{/�M�0�[
�!3VvZ�\œ�*+%�@
�&�oAZ$u��R�F}3ڄ[2��[���3�����ݹ�K�RZ��ȯ+��9�}�6ꕲ���+<Q�Q��&)�t���c�m�io���C�^hέK��7�f����3	��7�޽#T�!B?]��F��k��BK%�����1�zd���|�������W�F�m�*_�k��������_�	�
�7�m���8����O������>�U���F>?� tB��L]�fW$�|	t�g�  �<����Tf����ȥ�Z�ˌO�_L�4��
�O�������YW��<�xI��h+%$���5��B��`���BZ���ZکP���Q�u�gVa�$�B��!�W꓄�p��O/��A���x���֎�a����M�^�g�d�����+󅋏b
@���#�H��N�/4i�#'N��Gf�|�Wn�e�fT���<�I:�H�֩�U�+��n)�ZW����X�����aY=�@����rꗣ�|d;YG���@��@��u�hp�K.Yb�m���xh���RWOM�Z|.�)���3\�^A��+���6�0��EL_iT����l���%x��|0�$G0W�@`��HsbV�, g�,�\����"���'
=壻���-������r�#/���t�?�v��Qo yg�'(���1�lm�� ʊ=݃Ùv�^_�V�muU���IV�@�S�4�
p��~;٢���|��7�T�a=��ð{o��l���=���v���J>Z{$��KKW�*t��Wr&)zA&�i�k��=m;���>�m���W)�:�0KFDe����k������4^~�eXϥ��k`>*�����	v�Uj����a��
���2���j1[��*4�����]�Ӣ�
�.�D�k�"���M��4�Ϣ���&��p�yU��$��*;`�:�(5�I�g5Q���o�K�#�H�l�+��%Q�����/b���vsY�T�I�7�A��)��������)��k'�Z:���&[m����ּw����W�#���e�2��Dd�戋��B7=}��<�wT��n]����z�gɌI���`C�8k�����gƙ��Us�6|d�漖W��M$�	>��> �e��wP' ����X�d#�Y�T���ΌT��$������xz�[픢';��*9jf݀�ݏ�41ts+?��|��s�eW���=��=����Y�-�i�\����F(X䧹��=����ȡp�F�(3�h@x6�v��� �Qxx+6P0�?;����p��uX{=3���V~�g��S�X�aF��|�ɗ~�}�'	xK����B.=. ��7���p�b�w�g՚6��B�#h�6���F�.,߹�ƹ�Ncxp��~!hX�P�'����ϥ&�ė��-ՕWG���+'2V��d��hMF�fB�&e���|�
m��yOP�K2�se�@�L��Ƿ��'��\�㿒g4uO`����%}�~�ݽW�	�j��By:J��j�rhS�⑁ �8���Hd[�޼��tY�5����n��L�tC�V�{E�No	;р�kH�h�I���r�Bl�k�	��
�$'y�.O��f���Z7^���?�[�O�s6��2�9'`͏ߛ����U�������Y�n�zə��S6~��+DU�3� ���E�S���s5��o�3��ر�WP���)�_��st���������=�0���F����,����M��K7�4�vm�1M�Li�������ֺ�yj�Qی��/�U��������	���r�8��Z|=�y�)�6P�g��[��Kb�^v�	`�t�ki��È����z���&���I���
�A�'mp$l({b�y�6u�o�c'�a��]m���v�~`a̲S��pk�'��@�}}���c�{�X���^�r+�B#�.}��:�ӻ��ǹ1���O������G���¶��Fȼ8Ib�k&7��i�,1�J��b5�^�h�$��,J��_eXB-���3���_��L�d}�GX�v=np��ǡz�N �kN��5�?�����Kkv+�"���[!�K�G�L�<�X�S�����1�4G�&�R�^�ʎU�4k�|p�Ν���}��EY���q��E���]|x�獞=���`�&6t	�C����BCz�p�X�D���J�/�9�� P.��	���Rf��;����#���P����/��ӡs�E6>wS�m�p�l����y���˺
7�?Lq-�iX�G���5,�
�j�pN�6����,�C{֘��㐯����{w�>*��[�O���X�g�^:�tX,����T�Ր8:�� �L����)vw)����/�*l�&˱N����q���Ū�Di�ec�2�Mx��'"|���.T�'�DK��F&z2D}�g�P�*�R5�ag�V �$U���:>"޸tOK�)+�����6��*�@M<
�%p�C���D�������i ֞��O�Ӆ2�C�09�����6�э�R�"6��1y�,!m�������*F#����}�����%]܅̭���I��9�f!�G�0+���a��^yQh�4\��X齷t>�0c#[�f�����d�2�p����v��yi9�p�k�چ�����߅d�Wv-���U>�a����7�S��,\�6٘�*�C���ż��	�rZ���5}���1�&�Hw��0� w;�6ZlIVy���|���m���V�qV���aa�am�B&F�L�P4���am��|��PH�<X��|#��Md�Ҟ��=�y^����ۛ��s���2�T�;u'����wTB3v� W��r|&M���M��.z�
�=j�!�z��YZ{�y?$;�Hf�ZE ���S�O�L�%"��@��o+o�����y�M�����5�+���e`�C݉�ЬXO���WZ� �l+��z�9�O��?y���O�(Q��w�"}�8C�����*�i�*���5���m쵷�}�+�8��h��M�v��y�u�P\���if]�:v[�����*��,'L�Z��;v���߮���g`[�KZ�s����~�c`]�`;�H)Af�N`�E�ޟ��}ޝ��gx$�]�oi�f	\�T�x��k���͎�/ �����uIr*g�ŉ�i�cV�g�F�Ԏs��Q�U�ʼ��y��+�V���p�_�m��[cD�/7�.X&�� ��GpCk�'��1�W�5�ԿX��I�3MV5�#O@��I�t�c>���C�z�S�43����ZqkT32�\_���[J$SD��dg����6䪍'6� ���`cU���T��E�Pi���d�,ڣ��o]� 'h}}	�F��(�ؤ�V3G@���rˡ�g��E�s$��݁v�5J��ɫ��y���4���;��>��� ���c�P��w�_�r�E�x��+�{�Y�ũk'
��q<Yj��	8��7/��9�mv�s���M9w��,$�o�u�`�����ɱ4=C��H�G���s �,>�^ݦ[ߙ�YĒ�}���LBS�r�fP�`Z��K��R�PƯ ��W���Ѽ�ʎ�Bq3'8�](����J��0��r><�=�
��;z��*�[����u`��ĀЙW�nZa�Ă��K�U����	�I0��7P�9I���T�b�F�ԝ�9�h�/w����/E$7�X�'iHٺmD}�����X�\�|�л(�ğ�ئa˸u�!e�qb-]\��"���:�xn���-	�rL(MA��U���$���������f�pq'T�s��ʛ�g$���H��� ���1[R��7�x>�2��"r�Q�|1��1L���@,B�B���3���iZC~��O2�=Xl5|~� 'm�2nh5µހ��Z��u@:�%�@��*t�bX���iS���:�.b�T�(&=[s�A�����ݢ���*K�=,��62�Y�]>��5�P�7�f��#�n[s34�ʌ X�L�j�-�P��o�s���ɟ˷�Z�����mж�8+
��;��q6�1s8�QRk�\
�'�/]��(������73���'�O�T��6{�d�N)+����,��������v�b!y"՚	�tȃ@+� �Q�n�Þ�A5c�
�A�Ɠ0AF�K���M�����82~y�.|�|���V#j8��>�(��_XiP��-��͂uT�/�x~(�^�_k�b�*�a屿�B��������cMe�Fɂ����R!�����	�LV�G�L�.f� �Ii����;���?pP����zX��/�� lf���oR<���
)�4�u�*��m>нpm��EO��k6M�H,���'�|?"�ebψ媾f�8�~�n��
��L,�����;���]
,�t�u�q�{�zc�S�7��r<8%�Y&+C�Xt��Մt?5������3�!��Oxv�Y���
��I�{���XZ�w"$��Nkߎl7hm���qٰ��L���wl��Ƞ����/ ��ͨt)���فv���+���c����Œ����`��k)�b�B�,�0���-2E���V����,���}��v,R~Јc.2�	���k5���>N���+>M[��<Ċ
��r�����B|���*w�cՌI �ƫ�,�������?F�&������tP�Wf����5+�Q�_4J0�\����`�j�{�~י�Ӣ�-NNLK#��N��us��r��:�ʶ��?ʞo�X];�@�&�L�{���D}�&$q�V���#A�]3�J�ġ�����yd��a[V���ʲ���<a�<ni5�o�6$؟=�RƠ�!���\>P�O�\�r�w�
6�t��]$B��Y��m��X�)-3I��kl	,�!B���^�&�TS��Y��(�:��y"'K����%@$Rg���D|J"gD�j�s�]v�
x%D�s�6^�����	֛u�?\c�~P.�I�\a�0H�2{'d����R$��$xhtoΐ~��)󅀖e`�R�m�j^1������l�U�:̧��(Z~�)֑�ױ9�T��ي�0�{�:y� �[����i�c���0:�C��*�K�l����|�I�삥��:�'^!����b��.�s�%˪���r~m3I�!hPܛ5��C3|Yr���F��N%!�oL�v��A�-F
���N��ZkU�y=ָS?P���{$�;e�j�_�Q%���_����8�K�ˡY9�|�~>�OO��:�pj�����
�9f���@\�Pq*4�~��H�)�rD�m�kY����>����� �le��y»����o�Ch*��	�������;T�mj�\b_��
�'I4����O锫���V����@x�aN[&|��B^��?tG���_1E�ʉ��(뭧Sr���MO/�X������c��	P3�i��DBJ5.�JA�Q�n��Ռ��A�O�f�?L����0a�Q��뷆?�k5�$��������A�b�P�7L��Z����*����w��:��� ��d%��&^�[�_��2��Q�;@%mN���Ãtk#�X���"����[V�}����/^����Mʹ2����"cЈ���#@C,�m ~���033�s��������[i���_-�}����4�����L+)
��^;2��Ҭbs������	����y�U���uIH�� q�+��6a��-����)tP"M�0���]�X�μ�h#}�gv�Q�2�	d3��2���Q5�*�i���:�?p-�e$�;b`�V�ǥ�NE�.��y��@��>Xw�}����>ULw��/zFD�f�.�̵����{���U�����w'��(�u��G�{��G��R"���|$�\^NV�R������:b�ާ�}�o9�&�b�V`��u'�X1�˹���:*3����G���ͺ]9��,;X�`���.�^�Ii�:�*7����f�U������_�9
��Zl���GX��G�0�'�\f�_N�6�A�Y��]L5��%p��U��x� ���o���K�4H��{�-c?XV�;�O��W�6�8����;�0���E.c��M�H0���?����������T�����Yȅ���Pr����	0�k��p_�D/4"h||Yn���M�S���#�%kL�_��ap\���+סb�$_8��8�\���,9|��.B��~(�(��`�ޖ0���4f�?��	Ϯh�ʳ���FA����zv�m��T��]��:��lh����:Sm+	2ԧC�<܅G�GY�vj�-���t����le0K<P�q-�RkJCh��:S��O�íi�\�شP��K��$��n��Ɩ=Ԡ7��[{$S`���R.�C},̴�HW�����m:����&�8�9��K��W��P���~��kxwZ�����ډW�������*S�@<e)�R2b}W�$_���7}�u&�$]�M��9�V��:�|0�s�1(4�8�}�<�kI�3���R��2��B�L�E�j�wy�`}!���T��_�͊��<w��� �.�k���r6i_���&1;�{�������n��v	�TZ�ؓ��5J���c�*�CgFÝO:w ��}!��f���yǡ�k���\�b.���'������A�b=�Z#ے�j�Ɖ2��k�?�R��ͭy��WN�h����Z�hmh�x���f�NEZFI0��ۧI*Q��h(Q���wHZ����R�@;��\>]�(fI�_�3��Dr6����x�@�������<2ڡ��N#Gh\�f
2�����P������ B�Z����u>�ޑ&�[���8@Ϲr�a�M��w������vX�{2�_�z��' �_�l4ݑ���z9ʥq�2�
�G~X�Qj��)���'*6��L_x�_Cx�.9<�$�i_Ji���.q9�w�C��(�qb����	4���i�����������[�u#1�vE���b|�����E�3��Ko��7V�q0�O��XY���6���d���v�����(��?��
o[��R�1ĕ:�=تt:���X����'�n��^���m���f/ν��3�������I�1��d*��$8�����Ѷ�{���el li�Ec�H<�ǰ9�pE�RJ	A,V*�����V����O��V(�;F+L>%�;�(�@6�0�T�~�@&;8��6']��&j�z��%����[8�4e��"�t�r�A��g7T��R@@k=�\��Q�-�2�?�U�����i>��x���N��sӈ�K���懡۠C��}��Z���Gl�&�7^C���k�Hs��9�qzq��[��|J�� +.�|���q|;����'�H�&a�[���̵����,���# �qs$�` ��c�%6��R��^�4@���0���Z	|�s�qc!�dՃ�è|�&��tN:��#Im�sY�Ɲ
ik�Z��&z���xީ�?�T	e���Ԅ���C���KhƆ�J|��Ff�܌lC1C�	"+����:yA�,<�h���vq�%ؖ���;r��~�/�49�a$Ɲźv� ��\VT��%�F*W�Yt�>���*!���EӒ��u�_�^2j]�>d%R�Rq�!��rp�R��T�C��6�|}�k�{�Ks��)�~Pj`����#._�8<��fxh~��[;�.���&G�5Ndy~��x��I=C^�f�)��)�r�'U��+Cv��������3u�;����(�V�2�$5]֭+�K�ގ�'���XS�~�$�Z�,����v��JP�y�?o�����b����-ʿ�4����h��%�Ǝ�xqò��@d�P>~S���\u������{�6n�V��&�1tA�"U|G3'�&o��Ru5��{���/��c�C�c���5�I�1��z	�?���T,,3���Km����T�7��,�pK��Xp��f1�[��`����q�$_;\����dc�q��Ev��Ėk�݋1�p��P:	u3����|�o
����3(�op���\��%��!w�Dɪ�����S��n�u�R��i
k׋��çE�v
{)D���y�{%F8^�!o����D�Wv��`2�������*�.ز:��o�T�ш�D|��[Rd� y�[��x��)p��yW�&uH��S�����'R $D{���1ć�1C���p�\	,L�S���h_0uQ���+}���D�/}�lE�z�"�<Q�^���u8�s.K�]�#d}�L�D��@�|�p���d�z�2O�[�g��{z�uCtԳ�z8h.���tU��F!蔥�+eUj�=f��lAv ����6���*��JHh
MRk�E_C,w֝�).t~��`^�G&�͉4�g�]D¡��L���f�Q�!�ǩ�(bi�`θNbK��Ì��s�(�q[�8EЭ�eV�&���O�'���/�72V���	��K�C.���x�Ԗ+|��y�y?�� q���7��aTb!�bX_P68���Q����!�+���QiZ��s��t'Τ=h�`��P�v.��_FbR�y��B<�aE��>�4��x�q/P~&IVb��ز���z�d���~�A=�vΆ�Mh��r�U�)��d�.lK$B�P�9�B� h���6���O�Ku��RPm'@N�U�n<��&l�Y�{���A�_+�ơ?y�U������C)Fv�n�G�sM�Ǡ׹R<> �O��+��>���4�I����\L>Mk�["Xx���}$@�ս�5]����~��p˪y��7!�S�����нX���t�?��2�B�LFT�&!{M�wN�X?6�sAL�,�<>�j���ϼ��r1��Yl����ܐ�X�Ϝ%����+҇����À�1'����$#���5�E�_��r( P��Zz��Ư��M�9��-��C���\x؅�nv�nK�&��`-DL\\ȹl4W'A�sE�;�UL�#�>�"��6�)���P]�>�
�1%���z�i�������6$�j�x�[�0�3� Ĉ{�GU� k<�[�NVG�}�����Sy�g�y���%�%s���F9��A��i�O�\<,Z�uU.��k�RO���`A�ʎ�.d�����5I����@٠z{�66�M���O\�Ϸ��.v�g�Ե���j�D�z��τC�Xbd����@����^|�jy���2��͎f'/�۾u�.Cu'��{E�O��H�yC$E��	(ĐL�|�_rwa�e����"�+Z�ӗJ.>h�����7���=����Y�R_��x�F�s���w�\"�(�����Ob�� v�C~�N�ns|MWZ,PP?�bt.�8}l*t73�4 1��Ӟ	6�V�SZH+��x;ߍk�7zHQ$G��>��}(�`��J��ț�O�Im���������AC}�X콊`�@�ހ
x~�G��tٔ)�q�D�BA��Bv�Z��&7�cJTlD�%b���ո@A免u�(�f�ߙ�zͦճ��O�O�r�[���+��	Vƣ�10"�"�u�C�H$�j�VE;س>ڤ��e��q/X�#�E��X~RS�N�n��&�Oh�m��#AV��Oǅz\�)D�X��
^+h�J�M��[�D�ŷ�ܭ�Ȭ��^�ٍx�+jZwDa�8e���n���x��i�M�-S��|�ļ��W��s�����J����Q�do2C !O�����\<t�%hX}��� ����|�9S��gN�3�O�5�sLIp��ʑ$����)�+s�a��rM'a�q�Xt��@��ʊ_w"�lKn'�и�I;�R3+��I�?�e�*`�D+��s�JI	���	3�W�g�>�?)*��҉��uE��X�������vRZ.��u�>}�10UR-�Cb�9�si��9��v�GQ�ɔ�U	���UX#]}!���M��V'�vO"��Bi0�Ak�r�\����8�b=LT���8~����Jr�<ViR���D�yT�����q��s��i��m�N`=;0�/�R�h!��k��ֶ�ަ~gw�bɶ��f���LJ�0�"p�Ua�p𔊧�"�1C��]�#��!9�>/�~��vOw�9v\��Kjʳ��5�|��?P{rY��5�F�����D�h�~ZQⅨϯ�]Y�f�q'�㙟R��Z���Zj�oy���V�~-�1#򀼚AO�d�n�Q�6�N�b}A��K�֜h���pS�⨤Xj� F�Ѕ|$�,=S�&^�
��F��`���yg��i�j���%�qw�2�l�\?[�(�������2|��ҵ:쯂<V�%�8�{B�SЯ���=�Mƌ� ��*��~��K�3�J�3�U.��H/��S �5�Q5]@�����r�ej%�K����/o7o�~8�a�)r��!c/��ea�m.�
~*@�kgO/��Х:�ɖ b��J0$��"����h�o����v*��>I6aY�T�� �{�3�L��0i�C�o��)
�P����.��@�Fj��q~^6r��Q����$�%b$N8-��n6z�\��J�r_aw%���~���p����u]���%�m�?4� �M#sF�_��-p� :����:)N[�>G�~��Y��7�A�I�}��?�G\���9����k�|
/��>���E�Q�$�<tr�n�>�H
X�-3�'F��hWͰs=\���O3������
Li�9acAJ�2.�AWFt��`֯yO�0[��I�F��Z�RH,�]o������~�3��^�T*��ww*<t`l����W~�]�����ߓQ�>{����+z���Ni�M�}n�ǔ���`�&�9�j�F#�hՑEv��ua����i W ��H"�|�߲����<�'n���ӏNj[�I���2��cK$��-v��9��8Dˢ+��x���S8����^$H�D����V `TT�Ȥ�I��K�g�V��a�[���cՄ�2�!��O��uZz�l�qj��2h��E��E� /�p����P�	dX
�ԏz����������);�����I,�	ԭ��^�@[���� !H?["���kj3�T�$����]ͼ�B5�x�5nߑ��wf��i2���[7Efϒ>L�Y'���؛���nȻs'T� Tr~ԯ*=�����{����0�}��׬WJ��aB�W3Jv��7&�3`n&p6��Tg���D��UF�r��\�5�����:�����ɏx)��7�p/�~�Ц�/.V0������Ƭ�Q������U�h� �E�.z^[|�t�(9�$y�p�N��Sv����[c�_���\l쳑��X;j�.<����~W�����;�z�����ٶ��N�L���X֬�cA�LB�C�Ks��%���F|�9���8;p��*��/��V��	�PF�u@�>�~����_�:+׷MN
6�˰�9�ό�7�ܨ}
��k摥>�{�<	�����}SK��û�]\+�o�G冀��G����D��W2���h�-�$xu�$N`��PG��c�r}"�G����^�m\��i+G\ȶʒ�}��Oׄ^���:��d��s>Z��B��F �2�����b�H��XuP�8�s�B-u��@��%��t�=��ӂ��[nym�8���+�� VÄ�֓�}�;�_�����1>tB�W�&�?c�����Q�O��V@lX�?��})���!y;��xd�4��Pi�H���.��I[�*��pf�]=0��I-?����M�Q����6]i�P�G��|�[? ʸ3�Fʃ���.�Q��>"n�0C��Y���C��%}��fm��t�zBȇPR��e��;OQj��w�۞pj&$�$����LO=�yyD���9S�>9�ܴ�V��-X�Ɋ�|}hjBJ0�K��l�>)|�oM��+I0����Sm��Ef�^L
As�Q%��t�CO{]�.�m59�����C��W�ts~6�� )��%:3�hX]�s��c�S��d!Kw	��8����G�x97\)��B&�^P���F<
F��I���k���f�5+���Y�z�	�څ;�Ub�x��p"��aoH������0�r����O�
6��w��sI&ݴS�Mǉʤ��H����	:�my�e$�D�ٺ��>&���I5�&z�&��"�_�"�`%6�SՇZ,l��E�@��`՟�{�[1~j�;���0֥E.�"4t��6�(�9;5������G-�Ntw�@����*��n�".�-t�ף�}nyD�KyAt@����S$&f!�\(4܈�~m{����d(������1�\�I"�a]��H �q�v�	mH5���o�1��m��n/LX�5�'�PgnJ��삋�cv-��?�����寯ˉ/G۬[E_F�Ⱑ�0���kdo4!~��GϠ��R��;�w�29�?w���ACY���aL_OdH��C>��T��C�F&$��ؕ�c9���d��`�;\�(Ā:q,�����\*p�L�#�>U 0��3]��p�t6P��_�1V����c��� M�n���Ŗ�r�w���+��ۡ�B�M" l��"6�V�R�t`e�آ�컽�1aJL�G����2%Rg���ϐХ<
%��E[{Z@ش@T�*]}G�nxT;���A�:-dZk�2
j��><\�W}�T[,��}����Y��	i���J��dD�t4}¹��_��ѻ-��9V�4�ſ>�+N��*Ј-��ڣ��,��������>��=�'i��Z�x0�L�L?v� ��u�P�/��Eçt>��)H90�]BjKF��=��P@[��3��e�#I;��)�	���$:[m;NX4�C*��Aa
\Y�!�XJ?��+��h�J���i���(v#�%���X\�^��=SL�'#\����z�������Pj�tr��V����o��ԇ��τ%��#s`�]w �$K%¤y�
�{БR��J]�ӟB��IQ�`����>��)�0����Jc������M'����Α1�C�#V2�E�!�\�+����u���0ū�9�	'hd��-������?-E�sN��'T#ѐ�/PD=_���1�<=)�c%f���S����V2�D�W������JV���S.*��Ǖ]w�x�Y����3}�ᅱo<�q,���.b���?zա&��Vf\w(5����$	�<�+ae�A�ȟ4��;.~c)���鍴^hV��lw��̼�/<��g{f�+�H�̛*�U��}������^��LG�m�,��/�])�_&G�\�&�.�E�1�΃3�ǆCn�P�kULiӖ/������>��"ܶV)r��G�d+�R�ڹ��������yF�Ww5�P���-�皩E�<����=x��v������P�ݣ����g��d@~���0c��d�l_$`�ɰ�h��b�e/_�� �,���P!���D˜p�ʯ�X��qi�C�AS�6l�]Z換��Qf ��J��I�}��2mk(plz��VFK+� ������e-�o���t�F��8�h�E�+i�P�l[���Rt08�[R+��ABIp��97�����-)�*˒�����uoe}U:��A9��CZ�oXfp�����@qQm�^�����e��<gBPꉺ��!)����0w'�q�ݓ�d����%+�6�cf�I5��̹�#EP���x2��-�e2�ja-0c�))����b	[������sS���-�)'�u}�L/\�<����y bu�X�1�u1a�$�!K�N�	����Ȍ)b_��P�2C��0�~U��
�#�/*�a����&g�kXH]W�TS��kP��'���w�z@��M��?��A�5��/I�(t���~E�TC�q�#��h���/����U\���������$��Ta����
kZݿ!�I��Y�JK����������Y0��\�|���\���Vrmh6��-���|m9N^�}( T{<" U��)�À6�(�~�GBA����h�YLjң0����݄ V�pq��B#o����nU��|�FE�r�J��A�a�B�I)��=�F'��R��?�Ǖ����*�S^-ؐ�@��xRT��D�����E4Iq'�T��d��Dtp�ѣW��>��R���{���}�u��f�u)̖�I�h��X�o�X��	�|�{�Д���<q�p� B{@�QC���.�-W�`֮N��b�6@`��,�#2�.ܟ���}�dj�ҷ3ބ��[���,w
�\!Md�󸖒Y���}��Tx"�]�T��c���l�ۧDۓ`?;L	�V@VU�7
(U��ޚ�^���G1�5�Z�Z�\!C�g<{�%�|�J�n{)i�z6/���w��/l��G��	�!j���ԝ̄��fה~�)J���+��3���D��l��
[�;��AH"����G�"��*�ωi/ܹ�>X�Щklһ�uVu�'���/g�@��G.�����{�?�C�Y={�|A�r�]�?_�u�/+�3����!���$���ʊ�d~�A��|���>)�&g��Tߴ�ᤓx�X�ݡ!Ĩ��u�sG�H�9T�7k�a>�?���k{w���@����d[.�.���������I�T^/�j�é����ERP@;����ݍă�!���XYJ���	�)~�"�f���*�^OH�L�I���-
�Hf�j��7=$��#��ä�
�nT�o�R;�Y?�����؎��I�Ȫ>���9�j1tެ=T w˯m�-�`�S87@tJ1?zu"�9D�~̒�����]3�}� ������S�ݔ����%�^$x���FL��_���6N��.+�d�<��}D/�L�����3��D���u(E�<^V e�8}�VQ�$�#��t�Xr|b���"��ԗQʔ��Q��!aϒ|�^���BC���N�I��k�P�hA�y��p���ﶰ;�SYG��ѿ�\�]�%ְ��O��Sz�/�͞L�-�������j͍��P���?�q�}Zh$�@��c�%Л��	�དྷKK��<7�;o�  ��V�V"�u?N��D�s�<Η���3\�\ӻ۬����n5���sȹ`�i~��}aES���w��}n�zt*M�m�~�Մ?����]�n�`���>�
><}��;������9S�%�>�e`H�?h��bk�{�p�o�`Pk������3%k����=u󖥝?���#~�t������k�����4�Mm�
�G'���Q���������KҶ/I�O��e
f����5�Sԫ_f�N/i��/�؈Ue���8���Xv]�b
`@�<��Ch���Vz1{Σʅ��7f�{:}�o�ti�#X��6���Ђz��^�nu*x��{К%!�&T[ur:p���s�%�	�q[�,\J>�$Yb�ù�T�Z֞�p"އ��p������S^�N��qn�n.>]�_��e���G����E�|8|_���P�]���**yi�M�RJ�5�0�<DW��{K%�M�SM� ױ�5��|X̠8@o/����$\Pn�>��;dȹ��埝l{ߔ�(;�jOқ !R� ���?@�#!D��X7Y���MR'!9��C86�{(�X�/R����d��:��'����9v���&sT��g
B�:a�;��Toe떉Q�.ri6��r�ԟCo��t��^���;���D-d������1/�Ў�?b����C��L�:n��rq����#�����G�o9u��\<342��[���̚��є~���OV��Y���J[�����t��{ K���h@x|��D���8օ������6��zI|c�!.�4�>�����t7�e� g�E=��*
G�t��[W��_~�dezI>c$��/���F���#�U�Q� ���G�Rw҄>lmK����gt~�Hq��qt�Eei��":g�>ѝ����:9��#Ծ36��t�	׀�n���.�w�F�]����k��V��{U��H�m�㓡��M�� ��	���9$�~�'X�"˓�-^$�V߬��Dr�^;"gڣW7%&>і�[W��2#:k7m�f�'x_2��=�6�*�`�N������Ӝ�&0�=������֪ΊȂ�#�#�"�-��ħ/�n��+���(�2!��\��U����p" ssz��IU���NPz�'��tQ&���+�c`�F�j*�)�b�@L� �P��Z�����𗭃� c�j���A�#��'.?q6���~���;��u.�����V��h�p�bs~8A�d����3�G�Q�z}�q��8
�^<����nE���:���E-���9�g%���R��`vM�� 2�5�R�"''�R��#��<	���$�k�O�`l��/U��&yIK�]8Mg�R��=��"���^����Ƣ8�|�2���x����yy���i�C&s-�W���x�5t� K��t�.��@��L�� ?��=R|Y놏rB�Z��Ӌq��{`���x���8�����<�P��K�.�
���\�1��*�"
���4+ ة)��#�����dX
��9�^�C6M�/��=~�P��F)�=�O=6�+\�xrx�#F鄙�k�Oq���LE0a��*�%���5�H���ݕ�+���a,@�kҨ���H�x���s��d��^,�q�q>1� a׊��⥀b�@�����Ü�Q���7�2���#/{o0\y��Ơ���Զl��D=��a'q$���	V���&N}oM�b�dN�����b�(����Jx���v�z���X�tS&��%�gT*��~ٳ�yl⁋h�N�x!Cd}�M*��B�M��������c� _jƪ+8Q�g(X�}[g5�y���C�}{[�E�G����b�Oh�HV��,�g���2�[J��*`{[����,��f����q�Ԍ4��L�18��u���`"=_�vԦ�!tW�&�B�Ϛ�5A��^j|�ƥy�B��_s�0X��p��F�K����\�%�{PuSQn�#I�R�h89�hI�����ը��)F��vݥ��;����]���C�怡��w]鍶�:c�7�w:I�A���+#/ �[�$���x-��U��p�.˾�p�,O���>| ��߻פA_U(�5�eS<��b������MR��q��E�]#A;S�2�jW��6<��@�$�6x�k���`N�ʯ�/�����^���X3��t�ŗw^�q쫙��͆�-DS>�6���������D7ôa�7�T���
���r����]-��O`r��/�N;���|�*���X%D�� Yz�H#�/�dшJ	<�EQ˛�����t����p��³���
5{�0���ʤ���p��M'E`��`7ѕO�W'�D��Z	
�A8�W-#uG~��|�0(x�`�j�ເ�e�3��:f4bz���D���FμOk��9�8��v��u�@�����ƒH�ҪJ���p�T�N#��Z%�}H�=�?�$�B��4D)�X������I2�f_���c~�P�!"���no]��#NR@kg,n0X�QQ��a�6VN^���>��G��Mܲ���85�:xM�������v�5������lO1ڬ�Ӌ|�'�����!*����"��8)���
pRC�f�c�j��r���c<����������G0��WRGZ�>�;�&�X�����:�\z񶄓Y�]�'p�	�:����!Y�ݙ��y�!��S�hn�a�~��N~��0y����
$����5��L�\�TgUco��ָ�����h˖��E��t�@�j7��������Y�d�[U�g�Yl�zY��uq�G ��H�̬�|�Tv��7$Α�.�/��v3?��pE��f�f���uHD55�s���:c;��|��R]m���p�����?E&��O��Y��oĹ��c�|X*P��9�%v*/�~��U��kǬ:�7�~��ҳ�=�=��E��b�NS �,XA�`����L��*�6�X���m�^m�$��J3���}(L\�Q��tcu2�}����g�4����� kdޥ;���B�R�X�a��0��W��>�w9���]��;g<W�O��pTN�{3�Xڧ	�<��𲬼R̤w��t ��~J5l�U���~��`L�I7�'����q%�iM�8���QQ��k��T�Rݔ�ĕ��H>��w�36W71Я2��'��q�H�۹k�9m!��M�i床��w�#c�E���1?)�u�'+���J������v�2�N 	˵��=�N�NVy�{D���,W�Bg:,�=�]��P�m��8�q�[v3�GV���%m^��٤=4/��H|�F��ܦ��/[v� ��`�޷�"] ]�SrFEgo�e2u����'<��A��Z�2�g�@ظ�j�B��}�p'�N6_ڭ邡tQ��j�F��Bh}`SY�N+r�l�Y/9���D���3�S3���8U_�]��-���q["�H�͢$���g:"�3CZ9*_Y,�\ zT�� d6 ��Dt��3g���|B �w2���|n[S�jP%j�#\�����=2ח�.�/����\´���֪��%O��R0���ː"�>xd`Y�:�E�>(��ЂW7Xw��� �9=�n�D+g��]�ġ		n܍�(`^-6�� j?�b�g�� �xSOe�D�"�Yl/�.����u�!;�5���* ���r�˞��T\Q<y�n������T�$�ؼ��0�8A�eGi\��,���{���f���Fy܈L�ͫ%�je���Y����#��]�w�a���+B����h_H�����wu��M�U}1W7WRvn�e&#�S����u̍����1�xuI�n������f�
%���@`���rP��ܕ��P��n��n�H%���niG�&����i�f��!�b{��sP�Av���$]n�-��V���]ج�LQ���5A,%�h�j�m�)#/s�-��������Vo��|��Ê��L����yώ����5�LJ˯~��j�����A�n$�{��1� �`�|*��h���}O�CG�J����P���Y$���VQҨ&٫�I˝Ph����V��Cޅ�����˱�B����%���}��G�OP��2�HP]Dv�t��6�`�c���U��������s��~��Q�ƀ�L%�W9?�Xf3$)�;}���nc��X�T�v2	���O���,��2j"b.�-�HM���8�2�����E��D-ظ&F�b�H�P�nqx�5�A����|[�"���
T� �W��p����3LW��~�R�� �B�*�/ӄ:�FZ�����]��ܥ|�6�u�����F�z�2����<d��ܘ^]FQ��]�ģ�%�#KZ�j�_�#��lZ��p�X�ڔx���>��~E��|����m�$������q��E#T~N~����˧�a�{��*m���4�6c�H&�(���%0�p[7�cR�"j�*��	KVg�Kp����C�	ܔl��)����=�>ǌ�(
��=�]qO�z�k�\�X������
�������sd#���%�Ƴ���C;�(ҳ��Š�!e��L�d#���W��4$Pyi�����׮�qU��ت�����Ӈ�cuكK��D�	��D-�pU�]�/�*�U-{�OU�b��x�x�$���P9����{?�Gr�*"�aP�J���O�"�].IuҀ�B�$H̱����׊���n�Q���&���ݢ��1v�[�|H)p� }�O�<1���m�_�]V���M��H�K�lSa�6���^�6q|��j�S4!U�̤���se�»a7\y�.|c	�p�z���{5�;�Y4�'�+��S�Z�}?IF~�>F S�M���B��l;\�{�x�<;�n��/�J8��&�
W��b�
�'ZX�ł���!�"�W;����j.���L�y pvrl�h���84����;���g��<<���P��A�� Ӽ<\���c}��4~�R��Deo�$>�ӑRw����>b��[l�G.���k9h<%�Hs���E֎n�6�6ky��O��3@�=�=���T�K�����{��ʶ��^��� ��A�ʻ�<]��r����4�\2�v�R�ڗ�4�R���yTj������H����x�f�Y�%���%Hװ��'~{�F��q�Rh�nK�|�AR�8U5"���Y��G��~�j��~���B>�M�>�4�d��������)����d��6��+#���e�>�H	�J��S��LiAi�d*C+`_�W�F����
;��n&�4�g�iOJl�[]U�e�Փ%p���i�`n�k�O89,E7/'�6<�E�<^s�����g[5��%Yv�����0��_�.��"JI�\��9����*�ik�3~����;�qdҬpC�g� ����"͌씟�@,�J�b�َ���G��n"o��\|���6���uz��%�
7	�F��$�����?��կ�G�WO�DK��DRc�17W���[>��\���u;��'J�k�7ң�N��\��f��stJ8p�Ů��1!3�h���D����i#tu��'���Š���Y�b���u�w���=u>0�T�
�RR��滕	�����ӗ�+*&�a>(�����jVx�3M�l�J�%_�z56�ʠ��XҔ 7ߵ͊R5&�?��,�}3�I�Rw�&>�v� =D�Q��ٱ����0�
�U���!O�jl#a5�g@F<�pԽ��٤/�zi��Ĭ �P|����HX���U��5�h=#ڙI�e@�wI����`#������I�FD
��VՒ6�EX�' �熹A��� A|ޫ��mb[E�)	��h:��~	J6��TP��#�/y�RĴ��xQ�DfP��`�n��h�������s~���<��(!5�N]�ܧ)h0.ݘ�52ѽ�jz���FD��m���a��	6m�m;9�?�Dh �\k�9v`-K�Ӊt&��L��S<�Ϳ�dɩ���N�t���:C�x�Ϋ�o� "luc\ ���'�01؃ai+�Bݐ�L3ք>���=�~�p��_7w*l�a�|C���%VNA��yՀ�n)��8hZ鰆5�ࣄ� ��)z���n#����۳�Jr��֌�n����f�0�
��l�|oRk�B ��BP/4�S���V?�{��
:Nh��jH�U1>zK���������{F�9A�Ի� � յW��}��j3UQ_������ɵ�=�xCM���{���'v���9Nx���g�B�GQঊ�q�H	=�z����?�q�Ƞ3�a$Z˘Aj�=}=P��t��T������G������-~�� [���Z��U\��*�'f�,�� �}^ ���E�rH�2$X
w5�'����r�-�̷LƗCB̹6�].8�TU����vȽ&�jK�%��͠	E��	�SmI�#.�	�I�C��W�[���<��f2�h'��1��}()��K�B7������ۮM���I"[N�%4�}��R�������w0srS�Ǝ:��������G�U?���j��N�;�̗�,k@rp�<2�r�֜B�F䁿tI��m>�2�闈v(�V�~l���ϴ�'c�3��o��a��y�(ʜ�r�b|���h��/40̭5mnW<�8�SքT���&�qe[�:��!�9�o(w� �e����"p#,�P
/�J���#�by|��-��	K�ҝO��)��ų�O���>���-�d��E��T�[�t��G&�J�ji$�y��c�{�JqaL�r�CMB'� ��= �$�NU����G�t<k�đh\r�Y&�Dޢl�����,�k|�B��Y�gS��@Ĺ�t<�X=m/X׬~�U�7�wlKM֞�Ҿ�P�	�{L�d|��-/�h�I�q>퍱�$A0��	R(bM����Ǖ9�����`�L���[�:a��b1 �^�YeM����?�X�� ���8�ێ����F6_�����_�J\�Ր��:�z�$�O���L1�D�}��*?Z�p��]lG�ڏA��6����,RI��_�ܹ��%4#���Q�w ���1ax�г����+��T۠�#(v�p���Z�������?��N8p�GR8�ǂ4-D8/9V���&w�_�+���\�������;W%6qm�N��.�� ��X%���la����v�q�1vU������kNiS�E��`�������U�>������9�[j^��c���;�Q�N��*�k{�U�z�m�#���7�����U�N��xm{���n5��2�k߹�>���BKs�hO0f��a��O�kd,�쨪	W>��w�Y+wW���{ZS��&ҝ2�y	��f�rei,X��fz	�{h��.ׇc��(��� s8;5�v�%-��S�k�aңw"q�"O���Od4��}��8$I�IE��j�I�,��8��0Y��=��g); {'hFL(�Jaf�u��}�,3�!0�ռ��#�6�;@��ǘdY�9��N���`h�M��+�e�R��c��DA���p�
��d.���e�z`|��2M��N1�����G��
�j�K��6�")�Z%�C�eZ��fE ˜��p�/�u�2��{�
[����r}z�u����2�p�7£ ���4�ևa�D��&Ǳ*m��l�4*8~��
#-���R��A�A��췼����ծ�hU@ٶI�;�C�3������i'ھ������`�F���)��z�#8$=�k ���K@�B�p)�b����?ׁKOE�n�K�!qޯ`� Cb;��؋`�+vN��O�&(���u�{����\�/����)S��^g�V���e(E�;%�ʖ;:��� FA:���QRW߄�5;�2�ǍfO���҉��.�:�P����)亍�u8å-�('ߍܷD�k&������I�O�a��UȪ�1.TxǕ�w1���H?GC�5�T��Q��\J�@��՛1���h����}��C�r>�08�H�P�	�Ȅ���EC�Zw���
��Ïr�Z�n�'��������@L��fW��y��A�D�v�>�x"���S��1��V�b��Z�;�1�l��aE�:��������ki�v��.������w���y�r����_)�
��<T�[-̥J|p��}T	�[y=��L���[&{,3\��4r��I���(�4z�y;��xc�v���vW�*�S�h�s��`�\�`��(	�͝�R;Y��h �o��R��������d�|6�`?z*���*�=�lP�wʊ
;�U�빕����?)aQL�M��_r��f@��p��4����nV�a�4&�o|����4`2�Eԡ�{�Ayɉ�QL�c.���(x���y|D{>��eHV�LbM��ϸF	�E��+�W?��ZiQ��3��&�iA��*p��V��\桄%`$���;CC+o=�gJ�\ց{��Ǐ5v�]h �U�9�hP�Y��ւ�RA����aB�71��* ��,J-v����ʍD�����{���&p�bE���һ0������ ��m�m�rK.\�K���o8֒���H�/������S�M�B�|m��L�n���e�sg��_ϳ�&�o˔Vɷ�7".�L�5��ۑ�@����[��.\~gɼ8}V%r�ޡR�E��?�#h+�����Q�ɛ��h��й
R��V\FU�/`�JS��*׷5��*`Y��ܢ�
�'�2^z2�u�,��.�62K�a��ߕ߉t�ُ'�p��HAˠ;3�鉨5���aF�8���nc���G����W0���|\�=M��L&U/�T~w�V�oM��1er�:��6�bѨn���z9K^J��r�	cN��ɽ}�6�P�0q�_�P,�(�T?�cG�%�Q`"[
��Tֱ�� ��E\�԰9C�,���T�@㸦���֓�(�rI}�U��ipۮ���Gk��r�w]�����l�l�g�G�N��ō��v������5{�����qp���	�3�%��p�«Ԉ$�@>�)���0�PR��wD�	A�y��?S���rf���}w#�.|�ܩ���O`m��ɼ�̕В�b!c���|(��J7�`[h�O�J�D\n��K�Rb�%��u�jr,�����y�$<��Vq������]ӲfyQ�R��f��lq�ؘNj��<�1	��O9�8��U=B�)96�w�p�.����q��H�
��Ftd�ԕ���᮵F/K�����Nz�Fe����c�1)�gW��&J1�*uR��{7�_�3��@z�~<*�!5$;��ʤ�n!Kw�lK��ƣ��<�P�7S�������׌���t�j��k@Y�����y`T ��ܩ}�nL
���v��Q�k5g�u� ���$P�l�eGD��H�vЮ�y�:Ť�<(�K{VNj�p��*���c����\aY6S�4)��!������
�&0:��Eo6m�%Y]���FwG�(_ʏ�-d�)�D<�c���g&�TΧEu���6s�,򱿻OYNK�d�b«��l��1N�7%���aOw[�l6���-�ildkg�%������C7�/7��L�2���~�%��X�Yx�m���0��ax�}�"u���u"�fWT�$�~:�\s�%F�'�4|��fX㛅:0WO�2p��r*� :�(��!�*m"�����u�i��oQSV�E��7�����
�6�sgM��Ξ�@-������/�,[{���P�mI:�ѳ�ϚME�!1��b0`�Vt�{З!�}#^����1�����ǖ�EM��3|�"YyOjAz���Ŗ�W�OG �lo���Z����$I8�n���3Wc�Z��n����4h���V61����.Cb=���b\Jps��n���o!��{��F�Xi��S��g1:�F���AJ�����z��D
���;j@��I�`Yϕ�n8��|I�qm�r��xc�j������}t�s�!�!5pD���Q�e��+<���&x�}�;��L���d� 3;J��y������K[,�k���(����(	t ��ɒ�´�X��ź+,�b�ެ�X�Yly��a/)�rŉ̿��J��ӜS�4�O��I�4i��I���5U�N�����h���M���A�˜'�����'ra�7X��9��>�VQ
6�Ƭ�S	'JQ�4��JX�($׈�k�G�luJ1��d��Y��t�7�BF�m[X��NK���,��ݕ��ID��o��6o�1�h'y��-���iEP��RQɱ ��@)`�,�6��W]"c�^LEi���UIY�I-C�u ]X,*�A��*?�x5w�9r���r��q��g�ᴦ)��R򖿨S�U�`'$gO�T��آcN f�h�3P ��$Z���ǼL.�ʹ>�~�<b������9�7ݧ-S�G��0ۈ�w��n�t��gck-��~��P��=6޿T)��:,2кfh6�9�O��#ٴ���0vӒ�^m�i,�ctt?�g�5:�e)�i���І��n^dJ�V-N� �:͂rv�%T�b/pl
����yM�Q�,;�gL�L�V��X&���B�g� ��NOV�p�Q�)�Vcn�GF�tXY�������q����7$�cv+��B��Ԁ�����83�}AN�������� h|5�T1��������2ZR���I�0����7�,��?�5�B�E�z�L�Zb�� ���Q��h�7�P[1�c�R��[�NN<�Ʉs<-y�0��'
6Y��:�e<:�s>uF�:v۠���aJo7N�`	,7@<���L�S"�n����Si��-����e�?6�n�Ȩ���-�Q=5_T���p�2�>��AV����9�=�B>��_�ix��l�w�u&d7ڗP��#&J=O������l�I��S�If�y�z��M��G��
9��O�]�*f�]�c�^�Z��H�Y��������h���"q��1m^0��p6��s�?Q�{���h.�%��2P�@,���p`� ���]�됴XJ#�8�	�s����z.%�?XW@$�?˨o���
r:j#�����mj�ą8�m ��C��`�Q�cf�P*b�~��R��Zd�0Q�'�0K)r=Zk�^�js/��BU7�%psq��Z.
ڵ3L�	���I����ɗ4�|�	~l8��av>#<ښ����j�ßs���05`��ے��o�
i�Ꮮ��t�l��u��,"f�/�4i���t�l�U��16����^M��Q.�z���A�,m5K� ��vW����#Gd��D��U���"�1�� !;�#%�I��O$�y��4�
�| j�����%��Uҗ蘉p;����Vte��� 4��B)��݄�M��߼e@�@��D��Q[Z�H��]�k`���^��r�ת��� �F�?=��Χ�Ɗih����;()�S��{�t��93FӉ���`��e���f�7�ຑ�K/3�2l�>Y9C�%3�g�K��%Ú����/��܁��-q<.C&��s�Q���x'ռw�lD���._[=�B8���b��@���Z@pi+�Aː͝�����a8���<E��Ġ�2�q��![�ts�/�`B_����,��C�sl~ -��9ಋ�6̐�M��y?����}v�����y�$���F�
�yߏC�^ٵ�2l� ��r�I�On��_����WJI���'&��9�.�/s�q��,���p�m����y���������Sp���ҵWS�u�rO�Ym��pU����Si���b�r���U�z��br1�;v��-�"�Ib�;g�����V���X�Q�7�\V�n��'ܟ��\)j�C��i�Fc�c.��_ŗ47�y�l��sz@�3���B|�}v�`8Z��2t.�&�Phq����S���P�$��h����������B��dW˪
�x[V�3|�k��6{)��2K�`�J\eBw�@'U���ޛi���&&�0D8C}?�szԏ���a,�wb�}GΊ�ȗ���x�}Ҵ��=�m҆	���|��q*��\���֋۾����=uO�i���>��|�9j���[0�D�������^m0c_*>w*�e^f���PG�W[����g�#�����UE;z9��Ր�#iz����`
q�VT��_���0�d2�҂E+�����wQ\�"�+Wc��Q���>>1u� 1���,���vV��0`�I3��{��I��jƬf�)+t���n^vdz�b���i�3l�ɵ�m�LN��=ЯEy�Mx�(�;�U;���Vݵ���u�z{�s��	Ko=#���39Q��$ln��$�n�����j���t�Ǫ��Ӆt�Ѹ, ��{4p]0�"�X^c	:T�h�*��s�4���F��a�7Hh�=|�8�
0�_�ʥ��w��0<u�_����~�f�������������1�5I��n�@,�߼�X#/h���-b�7�܃�>zGWǺ
`rHZ��YUu8���[��sD���Vq�<c� 341���]'ʊN5�.:�x��@r*:��F�'�T�Y�8xߒL�v/��0�{�!��~�3�w/RMM��{"�#}�Vn`�:U�ÞTQSP��u�On�f������#k"����$��>-��?L�Yox�j��a�T�CŘohz�7�����@}�|+Z^�����Q���;ͳ�kU���l���Meωf��9[%�)�lAM�Ygn�8֛8���H��٭��J�Fl�~����u>$�FjTj����@D� ��T%��[���;+��v�ٵ��XTNX=�9��  D�s����Oc�}�^� Y�pLu`�şe����טF�P�[#IF�o�ь��f3�I��D�X��ꓱqg&�\�_�������a���F��c�Bm:�ۙ�`5��MI뾱c���(֊�һ��0�F*�S��Ƌ�0��� ;�B0�2��p�;�GuOs|��}G�������c� �_��y���*�� 1�>\�'&��J2�;B�4�b҉��Rc8��7��U����r9�K!��X���)X�?I����l��|��b�Pe��C[�,�fE9Z��[h%�Ƿ&�P撈��;%)�*?ڔ�"jC�T�qJ<�~�}{��~�4�:�|���u�UR/��_������̏��%�Lel��zDN#������w5ˈQ�m����A9�dW'�C�W��H���kU��[ҙ��Qrm�Db	����J+^��j���G,�ķ�L�>�����/��S�.*��L�!�$(�mC)kΒQ�ν�����p��ӫ������#Y�� �L�q��<�y��,JB�0nag1�7�$$Z����D�����ߨ�n��s���#���V?7��ԏ���+���^T�P���V;��$Fy�)D��9I#9}�|���l���n ��N�&�d|�G��s'����'j�@����ꐠ��'^G���
���.�˜���*����-*�Os����Zu�0F�Hܥc��,(�[h���ll�qW8��߁���9}q¡����;��c>���絲�A��*�UU���n�r��c�Q�7�AC��@e�@����sß��h��ǈfe���Uq���7
:;�qt���o.
����	����۸ŏ��h88+�2��͉o ^R�?�M9��b��e�D���v��9���52Kx\�?���9ݿ�q迦� U�	���5 4�����3Ѕ�-�r^pv����p����^<�N�L@[�MK��ԺJ:cp�*�u���>��Y�)�%�M����'���4�e�˄#�t-;N��q��&_�|Ti� �^;{���K��b�=C��QZ\�e�BJ9����b��d�z ��	�J��	�M�#xF�=4菬 ��B�Py�Uh����!��(����X̅ó�;�{�wEqg�Ȕ�.`�D��{�A�XZd��aD\ɪ��?\?��[�K��(,���O�^x*,)Q2Q|�����#Vy��4�^�2���e�ωb�E�ϟ���ӈ]2tq��I,�kb�X]��h�l�=�m���FvszUWV\z;�b8��6-��8�ݛ��:�v^H��2��E5:��h��#Fň3w�,��xn�]�'�=�>��I���^�y�j��[���wf�	�JC�g�YIvX��I��"@b����\�DG��#�c�f��W������{$��I!=i��X�<a��Ӝt��K�@�I��e���^Z�a����M^���w�s��S: �x�Klh],r�@!�ͺ��UH�5��@B���I���{D�*���Jyt��ͮqo��e��䂵��'ΐ��P��׺���œ)9����q��BvA�����q�?v|")w�?�����/c&��R����r�Wԩ�L���%�b0�I�x��k��/(N�66iKv�$b�K%�>���@]���*�H\���Zb!a�[����M�K힥�Bs�x��������qa�><kTI$H(�9i��͍yF�mt�oZR!�	�I��;s81p���@$*υ��. р��IvF~��Q䗓$���;�w�qeZ�N����<�U/���!��m�Y�,rm7�)�u%effD*k�O��zf n�%%2Ln���L���;�z?���R��C��3�Z����L\4�c)yTx�Γ#���ɶ���Zk�`4|2p�Dp�����V��+��{��TJ8�>4��yk�|���U�`?�c�X���Kj'��="yˠ����a����}ts�?�G�!���|R���Z�$����V	����+��#�>�׎��Ɍ�=i�7�1�:a�MR��������т�-� d�=��9����A���;����jac�H���y=	��O��Py'��x��Tcv�2�1ZyoH�m�Y����}Ug�~'<���m��j�6sW�i���Y�����
��z�G���@�=���/^p�nR&Vt�\:Q����{�d7#��)���vl��'���P��M�s]v�PdR�*���|:���T�c��F�X ]FL�)����|f͡'D�:'ϴ���0!Zf2��]���ح�\׵�<@�mp��T�	n�4�9�ov��,�E�F�������|�_���i����t~U�%�0���~Y�0[SYD'찲"��(�dvY��ӏ�͡M7��re��עlA���}��ÉC�)�Dd��ر�ʾ��#;��bGXxIg�X��*�4:_vOEl>��������0����?�Mƶ��?��Pw��� "Z"��.���8<�4]�;9ښƍfBv��h��&4V�������1�Ѻ�~h��t�N9xG-Dద���{a t��7E@)��3���B�Ήr�.�����;��w���;'���g�}�F�F�E�h}�Yk�Z)TpH�=�� �3����~����V�jvΕ���VG��
];RX)вD��JE:��4l���*u�-����A#���H��D8a�U�sT��\�� ��}M����\�YxKv5�6J����֟M�k��Y���L�	�`J��9�?U��j\�A�;]��]#�xM۩�Sn�^�e�� �/��=9�~CYxtY��$5��"���D8���td�WE:tE`�q��I$������2F1�}X�A����$mh�U3ԇp{�|f�/D��|��S��rY��y����@���l yE� ����A�#�/8*��B+��Y?�+�;���FnejH�z�2y�E��nt]F�RQ.�hv$���oiY-6��>'H]89U��H+] �hkdX9�m���N���Y�D���/vxe[�N������������R/6N��~��P(ל�����8�E��ĉ)�g��Z�8(Y����@�����F�P%��7*%�a��d��V�+VJP���u}�r�V�X�xP�ْ\��pT1���\�r���veK\�]�u���p�)�ј����:�Xx~���{C��z�ⱌ4���O�_P�iZ�P�ƪ^�=�����>ō�f�!e�ZS=�����𴯾 E�����0�o���R>@k�є̥iZZ�@a{|}�L�z��DC�t��m�Qg�gS�vtU�.��7A.�����5����
�"�UF���8DU\E(�U�/ҭCKs��� K��)�O>�K y��	6d�>�G������b�
GU�5��(	Cfr������q;�%m�a�p$W~��B��Ⱥ>���]j��>�=��7S��.6�
n���>��S�F� %�`�mp2�bFJ'�azF�͂_�(�,eC�\W����ř�%~S��u�����M����r[�^:䵑S��M�J&�[�xӲ������ ru� �6�D:;Ä�A��� ��Bx�U�`�=�>@��ѿ�r�O�h�^���K8BV�$CK�־%O�
F�����eWċ�g���N���'���2��7�b�- l��Vh�������$���'�"�(ՙg���?���.�p.�U��I��nF�V�)�d�l"Q���G:�0A����3$�5���1L���,K����0����̄��q�GGzy�~����>/��w�ҪN��Z�i>0�����`�"]��_��whx�*�fnl;�r�T�h��/��K������-�TU�\� 9�w�;#UfSF��4�I#K	b~���Q�������?��Ը!���a!�o*�u��?�F��D��Ý������el���~�r�KS�z��ag��m�T�;�$�UG��/�6�^���9� }�7I�?f���u��~k[Gz<��~Bkq&�
x�����rgj��EV���������8��5�	8�+5��s�����"��o}٭���H�<��N?�T �jhi����d�MWɚ,hu$%�-��]גּ���6����?��F������u!Tq�ZSS���s+Cm��4��i��u���ś4uɘ�����̦��wb�4-��3��M+��c=VF��ytQ�dp9�jGPWm:�bM�}-�T�KY�j�(�ê�C��6Iu�ިo}��\��)"�����W����H��8C�xm,\�಑at�G�NxMh=	y���"ܦ۝ބ�H�L�o�m�����A�0|��FBi������u� �_�6�˛o��z�)�M{�څ|9D58����+�1��^�)����γH��{[?��d͞�pk�7K�L�ؒ�w��c�E{��:�@f.���W�BWɘe�����U�cوqYf"��-�[�����E����x��R���<��/B¾��}a*���]z�Zl5�2� ��J�F�b�3�;g��V|·?XW+�����B�w'���UQ�A�&�8)��J����Ώݞ�n����&=2�D���g�u�k�i}�6���z���ZG��np��* G�A�������T/�(�=�Ա�'b4LÐm�Rv7�������͒mbmxLO�^�FW�W����ԓ�@"7U�B����p���M:\��(΃č�����̨)��8.�te��yԈ�n��]�����Iu������m+j�U����A0�Oo�,���v)s�<��\�q��ͳ������^=��J��F���1�b~!�X���h��:�xC>�/|����K�&�nǄ�Pf���\�x�9��"�^�b�~m'��9G>���t9,S6�3M'!7�F�+i�(IN�
SA���a�1�r�"u([�鴝�+�+F�'FClݒҕ�c�*��*���#���w�r@�uюPP���'!|ѓonW�/Mb���]Jۿ�� ���T�s@?7S�z��f)��d����]���� �2e����8��eK1�&���6.�`�vu�"ZLu��=���چ�`�i�H��V:�0��Y6�gƃ�� 8�Wb(�8Ą��NA�4^�:�᣸3J �#Wڭ�g���V����1�sY��&�|�󶁷)��e���a��<��DG�o��4>����Է�g�X3�/H�׬� o6y⦼G�q�cHG�_>�Z�Ay.*���Z��i�FOF ���T�όU.,"�	*d`�)	���y�gۀR��/'�O�-�2���t�p�n7��`�N���)M$�&K�6א
�FY�N�<��5A=�a�!K���8c�m�X�-"��q�3�3�K�4���������I	�O��m�d��!�a�m�Z�I����]��Em�{��<7-P��s����m�	'j~�O�y� /��+�_b^P�^b�8�=�>�5%�&��w|�n8��:bP�[������[�g�d�m�U�&��=�U�<���z-h���[�/�`�fy�@X���,K�k����E�&�O�[���0���������"��z�?},���P C��7�n��]���mn݄�"��.gj\���U�/��p/�o/) _��!�'ͻ�O�Ȏ:-�($��+���H�器���Dj'��١�U,��w
��<�CJʯ&{��!�cY�K�n��!>�"A� ��٨�3�Q�����Kd0�D�V��Q!���H	�̀���s��*�&��o�S�K��|���	���]R��?5�(��J`�w���F��9�	�-�9�y�lB8m�����%��CiݽI�(���g�/�}� j�0�O��B�ܞK��J	�A��e����پ{�\�"���5'>���U=5DYj��*H)z�b�C��B������Y�$���G���0|2t^5�]�s!Ū� 0���r�gͭ��Ch	��cV,���1S���|���В��f%�a�1�Ƣp��X�ni��(]ya%�)?y��DV��or�&�pb�:i���k�e���'��6�I�l��*@��&�|QBՊ�Y�� ��_��"�7�/r���{k����2���<а�v�>�*���}�Ym����CHm~^�Z�ծ�x$���!�F������\�^�9�B�[�%��\��%����?�סF��)���V��#(3�KjKAĉ�z&C��J(�-B�J�G�q2�p�;��ض��6�����N��L�O�K� �!�E���n��m��|2�5���	vh�o��HN
ΰ,N�=s:՞h=�fyG�5�u�cI�����`� ��N�"������y�8 7I��*�ٮ��,�V\�T��',5��v�����~}	�-@�^���n�o�j�߭�oA�,�*Z���7���Ao����h�gTC�M�7�}��#fa���{Y�Ġ��fO�?�=���K�nSzy�*du�2x�����e�����;�&KޜFNfI��w�Cw��sɂW�A�a�l
�!�����d���^�9ޕE��̺r�-N���C84h4tf����n���>A�/hXV��8GJ;��~����$BF����P_m+l�0<f!�Y�>�G�齋�y⨝�YD����0Y�c���rٱCx�uI.>�M �6��L�;�����ߊ[t���Kdi���й5r�P����3�d.H+}Gu�@"�2[�{��{�}��F�N�t�Q+0�p�O�u3%�g���ծ�ȏ�"ؕ�5xh�����=k3�)��>F�&w��3�����j�����GFD�d�T�"9N������ٺ ��,k��U^���%�^~~g޺����d`�[Qb$�OϮF�}��H��o��vj���l7��v-�"h�*A�Э*'�f�9��Vy��|gZɂ���
^l؈kMV�gC��kd}T��躂�xL��F���@4��NǶ^t��!��ʉV��$W��0QԼ�h�5�M�Raf|Q����
X�[�v�i�4l�W�@�[���y�md�v�J���b)K��v;�B�4��Ðܯ�I�6�_X���?I�@hBij�����)�0�\|���J�;�F��@BĖ�"d�т�����7��}��;��m��bmj井�XFR#��.7�A@����h�κ$?���3�T��E@���z��v:CS��'K\+�`z��)��~��I��}�\XSZJ�Kި��H�é[�!_�E 4���`V8��̜�4�^�RJ�c(6��{�7:�#�	5��W���R.�z�Q2Dt�A!*Z���a����!*��ٷt�0�?�L>�Mׇ��pn�����R{�5�m�7����`#�(�6zWk��	�LX�����ј����b(�V�_z*g��H��T9�;�[���bA���-<�=�`搐,�z���Fq��̢�XT�7�j�P����w��e��L"D���*����J,���ؕ�h��Έg"G ������>3r*!6��}��q�-⬀41'k��?��x���&�x��2��v�����St�}��Z���g��+�-
唍 ��� ���hUW��Kc�I��؎>���M{h��D����sl�$&D,
�� BwGk�HF�33?'J긳�5~�_O��t#2�fO�u�^�7Z�0?�p��`y��R.�j�dT��]~>��S�?t0fW�R�<��򿷿+
�Ub�gۿXCX^H;%}��E��i>�)�LE��'���@��pC��M��KXa�1��f�-�q�̃�<��d��5w�$��
�����
�f_���8��_�����l2�M�,y碏�?�o�^�RgK\�I�D��i�?uI2�'�[�	z�d*���C��u��r� A��z�d��L�Yy���~�3�3��i�dq�Z��'�^���-\{��J��GD��7����{��~��oUX��qx�3�M�Җ�Ei� �tr�t�Q`���3�e3J>1�̭T��@���+r\�``5Ы��x4���C&��mva�HD��va���g�{�THgb�Iw�|�@M�I��bk;Y� ZMG>�\�e�oeX��!"���x��B��6�<6�n�Vװ��b
�[���+^�2d��)�6��GP�o9���D\�hٕ�+٧X�=�?>�}�u@�[�9 |�JDB�I�X�l�6���\���}Hh��� ����[AN�R"㺦�?��c>��g�n�ӧ�	�F��oő(�,3�f����-N�ZGqpBp�vb��uA�)����K,�'"6�Z*6G�Bz�]pZ�=��D	�ɓ�]Ŕ�
;@�i!��bGVM�?����iֹL}��G�yw��cpl�Fʊ���w�9&*)��2܃٭x��������Z��B�B�vV(�?5��4��8���ƾ����[�`����6��o���e�X|��3���`�֢���b�"ZTE���x*[�����U�E(��ŨB%���=����+5]t{mít�Z������i�ms���z.��</�,QН�i�$�x2ܺ�g����X��*��1�M�xm3wǡ�=��� ��3�s#��UD���������D��:棎Z��o��	�6�q�0�Y��N`9�m��n���ͬ��K���V�4�����ܜl�m� }���W%i�+�yԄ��� �F�O�e�{\�,@�9VH~b��I�B[�=� MxU��^|ESȔn�4��̉_���ѫ��`�d�-M}��v�ڼFL(�2�/G�(D-<�-�6�ED��׌9t��Ƀ�O���|]�ھDƠ�u���
jɠ��rU�&k	�C�l��r�h驮5Te*��|�Teg��`)�
����A�5������M��=���a6*���1J΅�}�J�TRf�*�gހ�;X�����mk��}ݮ��pu�I�&������˧Q>�p�EȌ�<3w��B���� )�����k�;\�٭uGDq�^��߈B^���}�Gz���(��τf���x���qo�ߏ��]{�<�M�@r�#n��|8#�1	�?'�5Yk����ݩ����n��� PM��c��d�������Wy�Q2���|��7�R���&���6]��v�G��Y9`�d}� UF�2Nn��0����^�l]��2�uÆ�f	"�=za{LS����R�]���h��\��J�]�cN�?�%v�.��Q$�מg�����e�<#ʜST�s����Hy�f�zv�^�7<����i5����:�� ����U��t�P��B�p>@�f��@_�%J���By���BNm���Â����z �.�������I$���� �@�@�:�9)X�-[*��1K?fC�Y������{�d�Q�|�� ��~�3Mǫ���z��"�_�OCE���7����h�8]��.�0�R|$   �q�4=�{�d��+8�>��|Eb}ǰ3�A��� 'b�Oh t�r"�����r�V��98_B;�ͯG'79��K�U���� o����o!K�s�Aʐ���~��>��E����)�n��iCw3~�zu��)�,Z�s��^�X�&N3ع_F�E}����:��bJ���ӆW�H5���T1�pE[ �� �Fq��)ܮh`����Kp��xv�� ,`�/�4�?���DJ�%�DS�M����`�@kMC�6���;�ُ�:/��"j�����F`�Z�.tT�VpY3;"����VV��t����3����Xy7���IWQ�fua�L�P���X\�'�^D�y2L�x���0q=S7-�e��la
��H��pV�N)2�CB�$H�׽*ix���Ud��gm��S5��X�,���h4�Mt| ��/cL���tn� �g��^,)8e,�FZ�Tu^;�ɘ�D	�A��z)<�y���<����`v�pn�9,��*]�4��-b1 ���O�kȨ�
�Z�PorR��l��đ4%/!'������^�<�6�ԩ�#�$k�+�"���f�5��'p_�fj;eK:�o�@�6E��}0��[�IT�]с�\��˪����4���`3�I��B!ʊ�p�����{ș��׆�zY���Xezvh��S�X5!�P����5�m��	ͻ�ş}�@|t��Nm%�#�k�xՎ%�c�@��%ST5����y��䖶��Ϥs��ك���c��S�Kz���YP}J�L̈́*��s���1J#����T�h���E�nB怟�Ղv�7x(�'�?��-p^G+1��-�)i�}�[�޲f�ZDsw�*�S����1�(�:�3f�a�	~�unȟ�&\6��ʮ�����|�Fj��`������?��W�L�W'�Cү��)����W}�QP��
AC�Sd*h��6�?�6[�V@ɷ�k�ԕh`��G�EYJ�R[,`�
��%O�������N���)�����5�����P�VHw��_��7�4�m[~.x��~��C���N�4V%)��!�y���y�&0��6��B@�w�Krz���23	i��x�ǘ�,7`E�-$�<'�M=�W��z���u�+N�<�	�Dmgx���w�����6FܩC�T �<��'��<qp�v��SB�x�?�G!(��w�#�c#Mt�5�;�����{��ơ�� �d2�4Ss�-��+�x��r#Y�o��N���w|s�%u�x7��CE�J{ig����@������c*�&�Yӓ�+X�����gSW1ĪEّBG��<Q�������F����h�|xK�#��蕪�!��T#�?�҂�3
�Wb��'���w�����wguw�oZ|*2�7	F��P���/$,���}�nD���'9N�S��אù���gςNo��l��p�a�3rD?cF�=�I�����X��NѽS�OH�w�2f��M,E	1��8$�/C�vdS�(�;�)^�Pk�V������X�\�RۘV��k�V+��.K�׮�U���G�����q[$��4=��$�c����0,Qƈ�a�c�U9�z���7;M
�����>�B��}߻�s�=��L*`��KS��Mm.}^�F���u����E��:��0����4����Xer���W6�^�i|��+=��I�(�bjE"%P������Q7}E�N_���>�)�M^Bo�&%}]||4GA�
e��M�Z�u7�Ǡ;3hpw���e��:g����bY�2�mJ'�L���O5�X}K�jmC?�ֵo�����0�Ns�E;Х��I�K#젩(*��[|��AԞ-jU�t�[�6��.r�puŦ�ҙ������mKN؍��P灃���G�9���6U4���>��KV�+�#;�@F���]����f�����s4/���`S4>�i�<��X��M%���	�x����AM �󄾅1�['�U:ǲP�YiTz��∦�����O�-�=ߧ 8�#y�1�y��I\��~��GV8bRHm���L$2����ج��a=ta��͸�(��t�o��H�yV
�(���O���ͱ#���?;/�7p��9��V�ٷ�99v>-����\^�`e%����FXLZ�c6��@Bؕ�˪H����̻�R�a�%���d>'l��֣E�z[7bg�ސ�B���J���9��/�9x��y^���s0V�����Rt1�/�z�qk��<�Bu�1�~Qa�Q�������ǲ%� C��	i�|Wv��@��3��Y��e)� C��\?T�M�t\�S�
C�o�a@�YJ�j?���wt�k�V@r��'�Ԛ��7Â�3�Q)��+ �l}��>z���"������:��Zp�1��Z���'��m�	`8-"�ڈ�kc��N�Br��Y���59���TIL���M��0E����$����)n9Lk��E`էk7��T���p֨�5�8{�ֽ�����y��&G��������p2���}k��49[׈��s����mm�N�6I@� �;v�|͈1(p�� �s��è��u2�Œ�V^[��� ���� �Uuen��8���
�[��wg�V9�מ�am-�?����e�ү9v��rpx�J�U춻���}�v�X���gN�����&O����b��}�P��"-2��퇤Jme�>߼�cӬM�̗w�HbZ��G�'���6���X�7����g���?����~:̸B�׈YΒ�1�q�(�u���d2"�MV%������D�zbM�3yG*�����lYDcg�g{`�дl� .{��30�"���]��ͤ�u��m�w�]����g�4�n���Q�����(��YvAT���B(�R�~ǀ���3���ޗw?�|�iݺ���i��TdAɖ�"'�-x ���ga�G@�*�к�E�V�kW�a>XD:�c087b4
XL翢y��� (�'�]w����)<|E�V����O,�*/P;ߌ�+���D&��.�иJj��Vm/o�ƹ��)@ʈ�B!�{?�i��d�X�&pK��V��Q�K�s�h��̼�=�`��i�DK�|� v�ܡ�?_P뵳,X@.NM�'��hZV���<��]��Q/z��WR��r��Ld������Ȯ�q�o��'�l�������Z1�����Ճ�$w�s��V��?y�e��@�bÚ�_�Pw"yܨ�x1��_SSk�<��DQtVB�b��mH��N!�2o�By�g�T΍���`�N��:NB*��=�ڌF2�u�5�B�a_��xc�Ѓ��;2 �,�T2��\�יr5���*��-X�]\�Y���0��[�`*cN⯣!ȝ�����lL�`U2'~�MO�L�d�D�*5�_eJ��P�N[�U�Z�
��? })��A*�<�tvA�\"�jH��C{��	��F��vڽ��pb�;��$J�|��1��g�y��9��_�}���v>m�`�,"�'��zKL�
:��ީ֛U&�ypǛM�oWY@MI���S����m� �9+��-b�.ev?57ۿ�6�u��x�H���o\���6k���nU=qY�t�A��.�8�*� e�G����m��ب���p�k�m� ��ȶ'���&b4�]�یG<���i41s�!��g�xz�X��%���r���D�%�%��Fva���H&��eF�7�￟�!�������76�Th��R�>�rA���?.�ť4��	E��v	�1�s��ȺM�F���/'���aib_e�����ox2�̧���gVA׼�ֿC��V)��A3��E�4Oܣ	U����C"N/j�}�)6&��M(��]�6eұ�W���!eI�Cp��И['�{nܗg/H��-`��J�B�Nw����Lz���M���u�Q<|�Dɺ�����0��tA忺4�w���<AL�!��L{�R�c�Y�z�0�hqqSm#�Rf>��Tȅ� �!��e(ݹh���_��/l�FĤ�P�L�Jġ�'4r+[�ʔX�q�<���W��Nǵ\��\�p����:��ȕ-��I��At���'k%~�ۀPlw��mw#+P�u�?��"���D��'��VU�I�MO�,X���zF�1�#�ҍ��i� �����d����vfH �-Հ��PE��V6��nz.!T���)��6�c�%�@�04���!��xܠ{�q��KA/yNׇO��<}�Z�Ik�ח Ƹ#�{DO�
��������#�#��+?K�OdB�U��w��_[�t�~���`���\�3�d!3���2��튀�Mɡ�]�*[��.c�I]y!�QNsh�H,C|� �9N�K�*Rp�@��F�����l�v�TU�>is��0	ڵ�{��@+��-r��8� ��e�t���8��?������;&?.	U�n!�k������ń��*�:��4��;L�~Xm^���6���d�PtM�̶@��'�����x2A�z�Y�?�d�#�dv�%�2pxDw��=��� ���Iy�t��)̛�S`��|n�l�v��{P"fp��\9j�F�h�!B��.�am9����z��[�a�0��i�W8i4ء�[`�]r�(�p$�{q=ķ�]m(LXjGɘ�B�!��R��WK��LbDPHi��}csu����7�gB�b3<��3�s։x1�r0�2ͣ� 	���I���Ԛ��Cpq�y˖j��N��%v�$̈́+C�A%N
>��*׶*|%i���+.xߐ�G|6�?���#�$�d�I�O���XL�D�R{��iR� ��1�*邊����< ^�^r�\�����k}A0��{�Y�P��2��b�9{U�[P�0���I�io��͏u�-T�Y���jgg��FVbF7i�mQD�]�9�	PN��4ID�D�
���,��k��N~K䧠�C-��Q�<F^=� ������q���O%}x����%#�P�u'.#d��<J�����~V0�P��FqR��ԟ*QRI׍�)�餜����30[��m�hz4��^�a��_��x��I�7��m�μ���6FzsF ð�:װ���qI*.M�X��;���	2*�]��G�����c]�������]g���T�8~Ŕ��@'��w���3��=h5s�j%N8��1��m���L���2�qx��&ko���1k�Ѫ�0AֆVz��o�n��h��@�N;��BK�ʐ2 `���<�eN��L��ㄐ^��|?|�.H���֕.<K4ک���V2??me��GU_E4�O�{@7�K�A��Ξ�Co] �DT����F�F�D���~���+*Fe6�NܲC�s�N�ɷ�q�$�%�X�ݐ&5f+ڞ�c A���1��ř��~k%�U��N������p�ZY��GrI��y"�$��N�<$�jB������=�k����e�ķ�H��
�^զ��HIۭ6QIlB�N?R[��:|׋�����i�_k��ۮ�2��+@;>oD6��� �k�٥B_��;�L9U*m�R���_�&�e��]D�[KI��-�Q�p+zg2۸�hl�H�#�v@�_�� ���E���o� ��耏����ձ��o����LwK��9����E��;9��Ș-X '��P��pOĳG$���!�%�QN��m+�z?��lsW���J���i�� �%�+�}m�V+�B��6��d%�7��)<j��y���� ����?:�w:CW�*�[x|�ѡ��O��\���9�{X^Pϵ����!2{��<LL�bײ �_t�ݵo�F a!"���&���e9�|b^)]�q����ԭ��y3�,�аJw&���f���'k��07X,j��k��x��xg �h#��׷���z��`X���;���/A��W��0��&<I7�����������[誧�?�kj��Nш�{D�оNu8P�S��f��H��䂺\f!���h~�@u28'eԽ'@��E�MI�NQ�z��j���V���^ۡr��$�q��+��w�V�	i�xT�o��֨�[?-�������poU�3~4��W5b�?=�»�F���B���hx��XH��_h�!J�a�7&��2R@q�����o0��9�s��G����S�y�y����-FP��!�MqB��<�
����da��L 7��?]���A���&�n����,��m��="��ųƶ�� ��q����r����.f�]i�K�P�<�g�Ğ(��QU�o�o���<�gq��	b�|5��?�5T�=b�J�<B|m^�C[�6�HP�HI#�4�8�mV+ߌE���s_k�x"��A��:��Ttd{q�����T}Yŷ.{�o�1wnp+�|#Q�j���ӌ	��h�8��+�/B3y*�*@�(E:�jPޔ)����.}��,��0Ʈ�֞�MM���<d΃��m��hY�̧��|�]��Q���
�˫j��H:��B�HT�� ��0BF)��`)�)dSg)�v�T(^QU� ����L�dj^�4���Z��o�?g�:=zڝ��.���Vxl�G�?kx��� ��#��#���Ӵ�������g��"�v�OO��M�}{Uܥ&����	�f��7�!>���q4���Tl������':V��s�^����IbVi��:�q��9�O���8�W���%��Հl����z�m��� V*���n��>)��e��8~r����ad��2�D,	�l��dY� �����Ш|��_��A����i���{�,��`++��u0�ċ��I-�W������	�T�u�21��u
��if2P����|y�_�-�����-�&�[�������_T$���vo_�0�˯-������|�"X��^ߊ�@ao���'�wXy���=�23Y4��]*Z���=���\=j=}1�5#R�M_�Y����K*��R�+�Ŗ�g}�p���&:�w�Ԑ�Bٟ�tT�-�n��>4Z/��u�(|��A�)/��mwzc����ei��P��C0zQ8��'�[��}<���@�?�E~��LqFD�:�B���+
� �c4��-��ӭ����l"��[r991��-�\�9 �#��wVd�p��ǧ��;�#`a?r�OO]P�Y�'*�ӵ�+q�?;{L0��X�ε�W��M-����i4�<�E�9�����ZQF���B�Eѽ�ѐ�,�Kǳm'=��_�݄�h?<��f@�Ji+�D^�j��)�h>�]} &�*L^ԶM�0f֪i��Pܨ��L��t�s}N_A�����:�ox��!��'%P7~.`��n�����n1�g���-�w	o�;w:��������#�<2��K��_bHOe>h�E��Fּ�n�y�� *����������H�O�BF�� >DB���1<�i�1[N�����ehi+F�Xe��(#i�JA�����2�/^�> cS�W�d�8�+����j׉'��1��!ڡlcD�F�Y���/RK���u"!����m ��_��J4�s��+}�������i��*�:_c%��ې�ce�JB5�^�zW6�D��Ŕ��:��
��`AV'j���/��q�j؛W0Ru���	|�E[|i��Y_��>N,t��\ױ��^���W9��劑����(���zc����NAĎ�vh�s*���,w�b��0>[ 2�J�j�d<U�����?��j�ď�^��Nk�`��	м��(8cf�����淚;��?;>
oR6Xl9��6�"i�*�\W,���vo������P0"�9֎;̈́2�i�t})��m	��X�}ţz@�-���a���I޾�kP�ʾ7��V�\ȸI����l<1
��K�)h�P��� ״�2��s�Z�����'>V���/�����%T��N�v]bf����8�.b�d��,�x�(���>
b�@���a����Os�P3�Q��\m`�%9Jc-�°
��tL!�Q�ޗ�u��Jו�6�d�?���>Kp�a�ˉHή�d�>�=�8���d��Tv�ߺ��6cu�=�sd\r3��mԁ�D�J[蛤�7�}
ȔR-�����/�c�˯Zb&�;3�&�E��[Ũ�~���RQ�Q�3��|��I=�b�Ҍ�a����1�!_�X�?����vrQǹ��̀�#Y�L*7��_�����k˦{��C �d��z�#i�ȭ
l�6񅸋dq��!�m��u����"��&w���͉1�Whsx�,�]�[x�#�b��x����qӏ�/Μ(t�B���^j�v��1XՈ��9�+c�� ��<{��9�pe;1!ڨS*}�ɍ۞H2ږ���ֹ�4�j	G��V!_��:���f�h1��V�}�z�������fev�%��SŤ�!jT�L/Ѷf
G��叶x;�� m��^n�O��Х0�ˈ I^hyB���$���C#ʾ+N8s�$�?"��dT|)N��C
�wX�օs�QΜC��6a�Ԛ�(���?���L3�_H#c�7xy������^'���H[������r�1�Y*�����Y����;Ŝ,C���!_s�;�^��~Ky���΀���V1���ri�(��N�����,#��|�Nmf�,1�z+l" ��� �y�ɮ�u3/��yL�
��J��|���X��h����|�UAB�Ig��~�R
/81pSX�wh�],�ͨKu�l��pp9�V%}V�;�fߨ:���Ox�rߨ	�e�p3Π�
%R�M�f$Y�L΅��2�>$
�	]�ɭ�x@��r�bG����V =�������li%V���<�J(�ܮ��ɿ��d�鍰Vh���n��sb��Iɐ�����Y���	ū	4(���:Ĥ	�rFҖсhN�[ڜ��ú�L�Q
0���Q�y~�K�Gx�	)�QY�2c�r��g����ػ��Nd�7B)H�+2|.�겷#?}���s�9�k!+E c�<5��t��<ζJ6~YY.O ��F ��n�����^���fC���s)�\]�d�����ً����D]�'ufׄ�;=� �/C��Nq!����6�J8�7J������j#�:�X}���[hhG�5[.�}|d巺�Ը)�Ë�ۋ�pi�����~�W,3����J�B���vF{|H+M*���4�?m)��z��T?�[d�Cz�g7�B�b��������Y���۹ȡ	:<��U�x�����}�V�g�@����̱�f@H����$��S*��͜��G�]�������D(l�@��AS��c����R�=l�����f��̣���t֮���p꩝���������G�r��oO ����I�o�^��s��� E5��4@�|Ѵ���E�2n��怲�KUË�b�������%��z�k���I���&���fz �Iu����F1���c���hd�L�r�G�"O��������khu釓�֎�ؗ�������	�@8�1Nz�8|�t2��J�,�kz�7@�״��@e���K�E걮�����%M ��o�	�fM��G�j`7w�� A�<�8@G�� ^�0�^ 3���&����?�/ ����d��Q�ͱM
Ww3�tg�a��Q��0�);��ǈ|��;��n��(u`M�AQ�z'��$+es��N�O�K�	�OT�&R�3�����)��sX�4�^4�؟F��0z�<5�2��D��&
�a�4"�:���Hi�g�\�x��;;IBQlZ��������?���T`��R(d`h�ޅa��]YVaw�̈��T�}{�\)���o���bh��%��Yԅht����:@�BvXIɁ^\$��<���9���	S��В8��q{�2Gp��]�}�r�s(��ƺ�Pt _jnک�n��xfF|���g/۲:�����=d��WA�~.�c��9�ޙB��"�T��%��T_�A|����H�4��%5K9��֎���K�-�]�c�U4^W����~���I�6����c�~�p$`�6.�q'�a8Tx(SK����uW�$WfD��1cX:����)Y	�P�Q*T��M��'��.�2y|�+C�mBJ�
��'ka Ǯ65���F]*l�8,��7�Mnv�J��P}d��;�>���.�&1�"�RU��NPgl��
�Q8���7W�ȵ�s܎����	iv<LīI�a֓�Ms����l��2 {�E������a[�3�ԕ�*�wA>������`���)dUf�_��n]��r��h\���i E�O�)ߢ�.�U�~݃��h�3t���mz���̜��]���RUӆ�y���T�7fKc?��h��zԝļ� K*34l��k=�~X9��=�Mi<0��hd1�ц~8e�c��1lFc�lNZ�U��9�LZZӠ��"���֊��H�-�]�����Rr�b5bx֖Bǽ��Sq�9�����&C\nR�{��ۀ�lY�d8�!���d�]8��1[!A,��]��+ӕ4XqdΠ�J�ޗB�֍�{�&!I,��&��2�.��Y,��8�j%�� [�G���6��#+FXkj�}���؈��t��xY�.}�Vh���ME���	�2���I�?D��}rS�i_�!�]�G[T�kC��R����aǇ~��m�e�ȟ9#��s��"0F:�o�
�dO�7��]�=y�5P�m�����ϲ�V���������]Im�,o&�,^z7�C���\��څ|��D�v㰣��7q����c������}��Kd�<�_��780Ov�$9M��#Q�L2LǗ�ըO�''��y��+�L��M.���ՒhVrČ��Y�F������C�u��ӻ�[���tx�8����;�ٮ^gA~cM�A���i�ۈN��B�N�ժf�_?�v_Y1@TU��_=�W[���_qn�Ȇ���S`����D!�w�ۘi�aF��ۉK�:uM��*~��$7����V�H�s�Gv$�1&��9u�c[m��#P�
��s�r�?
z���:�ˋT�D������S�zs�M ��� �&,���`,fg�J�!5��'Їc�_>MyI��M�׶ ����N���v��lv>� c?�}�X������c�R�}�|���J�4?��vNvK���6��NxA�!�/d����4Xf
6qM6�������Ak�g�L��)���N��3�K���j!k�8�����k���q"�"Ӊҹ�1-��y�ɂk2�H��T����(���."�
c&َgP��_��B;2H�"���H!Eʄ�ȕ�i��F�ӡcI	��M��bCʝ&�S�V�H���G�{,JX���zuy#��>6�ݾ���H7w����z@��(DӇ���S��=���.�5�+\��j+r��!��f����by�Ȥ���[=���*cƮZ�U��*���C�Uc�7�8H�{)�Z/��[΁V�ּ}�6����%KA�:�Q�a�`���+��c�X���ܼ���(o�/a^���S���c��V��J���BFb������$jh��a��o1O"�28�_!������lC�������:��ˮ	4�������w�e`�9%��Q/�O,�&႙1i�n�\戕ͬE�>p�S*��Vڶ� g��d�c����
����,V$oBpS� ���;��@�:��],�!z�(�w�ɡ�h���Jc�s�T�k7x�qI��Q�pϘ���\�-,��(NJGZN��D9��RBT�*xb?�g,\�L���R��^��(���RVOywM'�,C��� �k����'��¡�W(�K����5�گ5HC���ݩ]��-1)�!���~#	�8���EhZ ��G�
��r0�����߷/��n��x&#���d�N.(���b� �Q F[n�f���bOzCt�0v�X�"�����n��܀�!.&<���%�D\�X;rE���KZ~Ϯu��&h���������;��FJS<���$`}#.s2Q����f>xh��@��`vy�B���y�϶����l]����g�`zQ4�&X�{��Oob�D��VN�7�k2���aaO4��Wo^��D���bT�+Ӭ���B߳��k��?�%'�F���CķLY|?�:q0"���u��Se��\��4O�t\^}���^n���z��9/�9k�/_������m���ܼ���W�r���7:�0�5�SFT1I}E���y�.�.M�����4�$�5K��ӃzG<�92��$k�^2b8�/^R���O��pk
���Yg?xcFV�����P�'� ����|~��ڍeqPf&��,iDZU/��%j�AI�/�{�������>���g��K[��7�\C��T<-ZＴd�x��\�̈́�=����*X���z�5��=q�O�z��xyZ�M��-+1���D��y�&�D2NP�A���8r?�Ȟ��s�V=D��2 � ׏%�U���B�ԃ,�fI}�#w��~�J`�h+_�L"M��/�hPS5���6��K���&�`���&�w*�@,��p4��KN�����ɶj1�P�[�<���=�F��d����QE�-B9�N�#V�S��d�WSo���U����e�6׍!f��*� '^d�c�0h-�`��[ɋ�b�wْi���,�_��d(4�u�s���nd�_�D97q�_`οUQ���1�y ���=����'t��
���mo��U@KJ_��K��-����%��e?�"�x�
2(���������tX!�#+�o����I�|���&_%��a�2���.ޠ(�x ���G��jI
W�O~������"���&��['*����A��5g�#*#���6.�`fN~소�}Z�ɔ�]8�����ʖ�E,��.�G!�,����W���j£�k=�9�' Y�2�n�=iĺ���=� �l�G5#=Y�d��[,g�W��Pch:&I��a�X�W�9+��Þ��&S޵?��1h�Æu��x`)�����Lu^$7Y����;�~�g���is�5��JEeU2��O���t�������o��
�l
��[���9�ZR�R.���F8�C���+@��+��xUH!G��"�d�V���kz���/�����a�5o��������Q�-��~64�Fx���:2U�n���A��?4ב�G�@79�?P�ęO%,-���ko|�GŢō���}�OF$���-h��c���Ԯ��I��J�\��n�+�>	Y�"���H+%��ztiar3p����@��+��qc�%�j�p	�^c�#1�1d�����@㣞O3��Z=d�0��)R���S�T
����vӝ��*e�5Qv��زF;J��<��h=�44Q�:Rna"��+�
����jȃ���7��*Nאm�4�qbW���uq!��Ps�7$�=�#��Kʶ������+��v"����rMv,>��{2<��:rz�.�@Q<v�Ш
��Yf��k����M�cz0L�C��k�>T@��gr��p����S\�@4P���x�q����U[��r����f㭃;>�A� =��ܒ��� S�L�	���~G�F��W�6+� a��s�}��,@#�������3������� F����:�K@q����T7'?���P*��*�\]��Lټ+�k;�Gt��?"�Z�끰�O�flCuԚ�tu�V'��U�n�
��J�p�B�����\O�6r�ܧ��}�����#�!a&�="Lm�dO�嵛��/W�X�I��K��6�����
:�*^�?�,��j�pH�W�毘�>S�e*��%���(K�Mm�������֍wtU��yr��|R��~�?](����OR��`��BISi�M�\x��K�X��xY~�V*����e��i���{��y��ؤ5L���O I�0����K7Py�H 
k
v��ٴ�$l5�X.�g��p��%u��,��7��$t��J��`q7%�/�C��՚f�:�ĥ�e��fp�?>C�Ӊ~4�D\ȩ��4�3o8P�%/v��:�$3�H�_׮6[)p	+(�ٙ��t����8<%!�I&�Z�4�� lW�ꢌ���P��>H���(���v6;L���nI��3�Y�{m��b�v��h�謭�T���!g�:��2u<�wG).-|�n.���Q;QR��,Ad��g��u�����~R�V��Y�V(�����\,�#��̒y�M����Æ�B���+b�VZX�Ϫ�����h�At3�\t�P:�� �-�k9d��Y+j�ʗ!@�E��ƾ
|q�ENXr�%4Z�"�AY͔n�Zd6�@ׅ��|�Z��H�V�: ���Z�|���>��,g�BZ�V5=xK�?��sc� �����Lu��dH�p���@7Y�	�ܱf���T'�����ZM4iS!�ZU�{�t��md�9�����AX6V��f��fO���)!E^���܅Z�t�X"��^����36�e�3(:����Fݵd򿂤p1F>��D�1����;T�&/?v�Oq��,g������b쉟3e�O,�8�\�ѾWw�L�t,���9����j�Gl�q������X7�syU,�,�j�_���-YѰ��F�]�&�2�iq b��H��+��
X���x��6D{[j0
v����w��G*�
�]������e��F��8���š�>�rmune�j¬�z����X���t��e�rDs�����>\�κ�_e�DN�\RRË@�0z{Z6�Y��ƴ�p�ť��;�9�Ƥ��c���f�/z�IỔ�Q�N�]t���&��D=�h���LE[SF�sk�C��&��-���1.1{yk����2{�% ^�����v�����FCuញg����=�C�k[T�mx�A�>�e�i�s�# �ӜOMLS�Ą������\�{�W^g�@*?�5΁vF�2ְ�����+��W!��;��UJ�}:7:I����~�S8��A�v�Gb��N�������$]�-�����	�V�b^&��Z6j�����Ls���0���Y��n��<���'�I�T�vY�S�����O����#�B�e�b,~1©%:]�A� �
�CV)H�!N�y�c�5���|�7S�;P!T�6�.�Cv��@��Ԗ�N�
��z{U)8�)/'rq�)}�Z�|~�F������r�l���#��b���Ww�� �ֻڑ�Y�A5���������Ga��A�����řG��Τ1�;o�d�N��v.T�q�ML�D����(L*=7�HG_�,ſCd"��\�:#�4?���6l��^���Y�$nrk׾F�Hd�f)�[�*Z'�<B�1��^�4�#a@T��ez��R�����Rގ�N������z5xZ0�������U/W,�������Ǔ�}�'?Vx�I��]D�ք��I����+�oP�B~��FgL+r�l�P��I��M�ʜ͹����Cn|��G�pf�8�7��Z>0-Υ�̑m��_��k�����l����Z�'�\����G�x�?09U��
|�J�-G[Gy�(P��K�D�kiS��w�3#=Q ̇�8K%*ɴ���Tr}?=+�)���RC覌�J�`{�����şo���^4Ğ���ٖP�?R�u�T̨�cX�G�Z�/C�Ca���V��1iT:Ʉ^Îƭ
w�5�'�v�x�ϖ\I�\�sPꌨva-��� �ީ��Mø�S(���A��N��Sz��"QA]�
����'-�� p�i����h�LI2Pj ?70�gvBk-.6��3��
[~��{K�k�6Ã�M��s�nMQ��U�2F�����w�*�d�H�һc�چS�Fs��F`&�A��L-�M%\�G��|FI͵<loq:��?J-�<��|�;5����}&W�ĠJZR��������S�F�����j�2J�ҋ���uD������2���;*�MÔ�!�W���cht����i^���-?��U��q.)�^�쩥[{V��)H�}�4�	`t|(����?~��4o"����GT�i��k�V՚0gDA&��z"${	Ҿ�q�Y	�;q�3��m��J�:\�);�9��A)�J_���A>ΰJ�r���+��x�q���C��Q�w��3UTytz�ՍX!b1d����u��4������Q��:	�@��	�%�b������$Y��PG��l�����	�����|����f'n�~��'���J[X/�{,i�ݼ�`1�I���hQ��x���"�>!��X��j��L��e Q)���uFA=�)�n�O���`�ᙨy���#7�@d�d�v��Ú�	�jVɽ��O}�>���9\}R����D"Н����gf݊���k�:l�Fj��h=q�j����	��ӯs|k<�I��ӊ���G��HA���s2錅>�(��Z^��҂����H/Ċ@b�g��	5��
����%[լ�@R�/�� ��B�v�)9^����GW�{`"`=�H�2����m�a�zuR)_��[���nr�V�K���F�8�B��7ts���n؜jh±S��
J��iCK�G<�����x�W.��F��]�K~�:U�V�b<�S>��|�A��ՔN]��-�]�dm�V�""�5𺊴0��'i�X�N�;xm[Ne�ޭ0�`�怢��v�>E>pTz
!�� �-[;�ф��@�k�_����u�w/1��1���<3�p!��|�(�B�T~H�2�����K�sPfǮ(�T�K��VQ�1!�V��v,&���O��e�D"o�8�|���Yg	�R��{V`��
-ۇ���� !�
S}�c�&�/����<�̵xк�m�;Pj$>�e�\�I,z��c�G�>R�$�tu�h4h�qP�Xۿ G8�ߒ��ߖY�^N��g�ӹ4?� �͆���{jY	5��	:�譳�6@F����*���ej�ny< �y9ӌ?@1g+�6j�v%3K�r	�p<~8���LH�8x��A�����iRRr�B4�-�b^3�v[� `hX� �0s����qc��M��e�Uk�j��m6]5�N���7;:Đ9��e~e��j'+ito}�lr��/��O�����R�G���S�'�Hv�_��8%�}��Hl��{�t��q" pO^���d����쳪
X'�U�D����1̕��+�M�a&�c�����<���)U�:)7�v���x�d�~r
[��S:q�������l�����1��5�m�Y��� ��7�8G��E���4�'ri3��x�$
n*5&����f�1�nݙk��?h��,'��T�huB�%7�X޿\5H���Z�1�)��	,�ݎ�0"���o�)���l���87`FϿ�*���c���(l��s���j����P��HE��n�%���AI�pU8*u�� �ю�GG���r�-�A("g L)�F1`p�Ж����o�!��<��I��7��fD�t���(��1!T�y�by.ɥ��,�ȩ���n�ځ1�4FŌ'g��0&�����$+t;�L���(a���;����ލ05.TڣMخYS�~A)�,��L����?3����9���c��2��Hc��}�z�$Dؚ$I��d��:w)vw8R�T�(S�5���j\kQ8	a�齧c�2'��m����%����v7����:d�r yC^�NX�F)�1-!g����_�Ɉ�g��@����U�:�m	2��ʘҽ_��;�o12i&�V*	a��p��5MpjWm�m�: E`�>Χ-L�U��+��3������T^�@�CRݍ�(h�5a>7X�Hx�s.'B?eWp������M��ᨦ����G��/��ȹ��WVп�������^=1�'>��Z���(P���(Q���O��*�rU�� �ҡӌ�E���4��m����16�"I��#���
�Ѫ�G��q�깯�R��;��x4�ڌ�����S��ǃ��;���i����"��k,�䚎S��h��s=��RF�&�5Mg�9}���gV���Et�Fsj4PJ����p���Տ��kJb�^r_\�#y/�'� ��7���#R�eiBT�~:��2(����n2�9�i�Lv�{�r@SΞL��˥x"���z�c��A!�hR��U�1e)�a�9\�x���)�;��4�g�s1怊�Cn�8�fL}:�d�/�#��j$BXr)�3���y�"K��8�F�ݮ��ox\�+A?Pln@����#�q�E� #6�w����;q �9�	�q��(�=K��1����8�~Ft�QE��.ʍ��Y���-L�����J��R��!tc*yc2��q��k𑸲G¼�8'[�#���A��Y*�E��].��Դ7 ��?fϨ�`5�{�#��*�S->�@/��oK\��g�ҮO��R��.��l�qX�ž<�oP�|���'9Rk�V�_�S�Wm}#��� 6:X2b���z�o��$o�,�+���(�f����bc@�1�Ēc钷�� B����$9���A��Zsm��i.;��i}r�����5G�:H�ڵ"��������v[t��,$�{�*�+	�ˠBud}������q��� yJP�a_.��;
q�2�D5�1���f��1�<U�w�|6-�1�Q���ڞ��ߞ5��%&H⟩��JO	��ri)]`u���ѰZf8�d��DqD���+4��]̡#
�������U�Y6�b)(5���7�a��ܑ�([�ı�r���b�<��͐\4�9�]�zjö�}g�g�m�1��,ȭ���i�`)����J!�B�*��=����J:Y;�/��
:�F�Tls����0��'��B5�e��s�o���Jmy#-��Ě��SK
~�;������L���� q͚)Bb/2��#\X�D0��,\�Ð]�)�Cn'�k0ۗ��,:�-<�m��G�2~��E���"G,��fn����~/�K+z=�ݶ%"q��GԵ�X�^��?P���'yF����������Z������'�<-H�S�kU�_z�j
�������i2��>�����;r�rAU<-�?@��/��@I��~ �(�+O�bK�љj~aa�^��)S�u�,�GiU���f��1W�LUt��;$b��<-A�ibq�?Z��%�K�r@��:�#���ԕ4l�aV\��-�˂��P������ �F�	j`�|ል��R��2��l8"� N��#��F0�
2(,�p�	��10�IWHB�/�W���G�k�	���n����w��aɥV�}J��������¨��zH06��ov���j���r�+;��($Χ��
d�b&��OPf ���w��w*#�1���	.hi8��ڐ��g�$u4�=�t~�lU�/9s��1�O����Ni؈qR-sBȂR�	�����YKQ�"��H�9�:�o�X��v�Ix��p@GDN�/M�������
��7����4W�)P�s��|`��N���&UE���rv+��0������h"�]�����G���v���\�%'�IХ��/#-�s���4+d��\J�%�T���IS���Ig�X��'lY
܁�A%x>����Ҁ~�69�_\[��ʮ�ٗ���}Ӆ�P\"QW�l������^
��,J��R�Z��Fz����s�f+�
�b"�		 �h=��
�E��c	@����7[����t��f��vay���;G�;�<"���%inC���)�����b��;�y�f�C�T��&��&��+$IT
�R�ӊ��"��U�-�h�c�/��ձ����Xj�!4Pp�,��V)K����c��z�$$����-�U�f,��������9"k�	�s#ޓe�����#NP/���h�SS`	6���2R�g)��XQᎶ���KjܔJ��L�y���)/�zA�݊�*7l�:�����p��,�w�Cɻ���z?�I����mWxIku�B{��R���CnmN��V���8�����K{�@����}p��4��WjtKu�t�z�~�z�M�Ԉ"� ���
IA��q 44A� 캶�gQ҇�[L�!��m:�'�E{�6�0J��p�.�:�ߖ ���YF6U��R�]B��A.����& ����$��N��	n��Pd,��_~J�U8��R�$q��#�Q��ng��t���$n���[��0X�å%���N�e v2�n�k���V���d�%�7=K� ��W���A�V`�.�@�"�cS�G��D��v��˃�nF�k�03.o�z�]KJ��[6z����'�}�:�i�t�WAU����2'�U;��¹>�Iv�������Y���&,.���
.t�k��{ύDu8���¨x�6*ٵ�a?,�3�Z�s}E:�k5��Ƃ�s�؝���B:n�o�xU�mߝ�ټ��4��&�$$�*Jz���Hʊ1�_�O7��*�)�&W�d�P㉜����X *���0�S�Cc�ጴW��d%`��}�����;��*zF/���^�I&�����zk+����Tٚ�`��_$�2��8��iɽ��r�f�>��+ax4�7��X&���a��,���_�ΰ�C�H�z�Q���z�rOp���{~��*8�=?��Rٲ��;������5߾�<'ǆ�Z*�X���ŋ_�ȕ��PMO�h�Uϊ|���LB�i�T�!Y�BC�I>Eg�Sŋ�s�U��7Y^E�*���m!_]���_���F
�Hj�Z�}�b�e�CBXF�e?dP�;��aĩѻ媿_�$oGҌ������o�5&������8Q��I�[;ՀU��1r��H��NҳG�<
>H^D�ͳF��~Ϸ.,+K����6�St@�{�dxsa�X�y�Y#+��5���c;1��\?��D��r��WH{u�C�u��YM�2���(�c��B��t�vUm��L�,�{�S�ݕ�u���
��ƽd&��;p^�N�zԩ�}̤���f`{�q�@��CI����t^0�5�D���@d�h�z�c9�`�ڤ�^^nu��1�|Z ������yH>[��Sz�M������v�l�	�#V�s�@s7��\-@��D�`{�K�x�*��|��T~^J*J�1Oz���CF��.1�lYo�<(�jΛP��K�s�С��h����Hqp�a	�GH��&����j)�P|�i���t��m��� �j2MJ���J���ь3V����F<�.T=���>Gl��<M���=28u��;1�iD�	�s��F�:���e����M�NUV��?��"�p~F��15��7{,���+	�W�@;�ϙ��f0`ږ�7�ʃ�-ڬ���M��]�>&�X;����E�S��$��Oz
��Nl�6`�����U���7���XZ����(��6�r���)�4m�c"�3��x�ޖo��Hx��v<W�y��=��������������1�` �$\��ѭ������;	�����E@�r�@4�ʷ�*���z�=
a��1UI��sj0�Dh!ƯP(zŀl1Ǒ�R̚(��y��+S��6g�����-8�9�@����J���h���y�w�1u)�J��rN�U7�L�5�_��]P!@hz����	4��W�k���mn��Ət�_8��25g,�ע6�T3�Z1h��1���>�� /��!�
=��
8z��W�o���ػ{����Zh.������ԥ�_��b��!��B�B���8�J�ε��b6򾣼�7�.4,b�e~��bѢ�`�4E�z���a�T��.Bmo���m=X ��pP�f�<�!y�������H��7@V����܃�"�(�/e���"����#�����wB8ЅUw�vp�J���kczOT����,��2�����ϙ9�o+�_��ӿTg}�R��K�;�]S�̍�J}��c�����!K�{�*�63�����Ġ:����Ⰵ�1ǻӖT�!�5�����L�����P�gF��
���q5�'�^��X4�$c�ﵥ#>p�,3�^B+sݹG֊������^i̍�`��F6�C�:�0̆ɏ!��)-p�*^�>r�����4_�P,4ah�Y����5�H@7��:�����*WI��d8�yGpQ�8e�t�@��eGq�{;�')y����T/;�"�=S�@�5��^���!Ǧ'p�ao�c�2�� c�9^�f�/7��n�]��ruvG��\������=,��UY���&2sK�ލ]\'�wb7�j�=Kdַ������P�}���6�u/1�'�*�0���6P��rN�������6c�����5�:�gZ���A��4$m�� � ��;�1��CW*��M��� ���x,���}�/hEz�r;Y����\�r|&T-�Ӹ�ˡ<?�T���qk��u�5�F�h��0D��ڬ�NQt�FC7e{��S ���GS��}�)v���1�~�[:��
�A���g��<ٵv�����hgG��ڥ��#|!���Uc�.��� �O���y"��N���(��4�BS�y]C�t����C�]��U*�o�u���.�f��'F%�H|nz���2D�y1 �_��h��l)��`g�V���{#ֆ�����o������k_�8�*8V
��(i����ԅ����Ƃ{��V���Z��'��6�V�����ʫb{���4ܛt�j��a��kj���p�8��L+�Z����oU&���3l�d��AGsi��-��#]��ھ�$�^���A�\SC�xo�2%dU�G���W����4(���s����q�]ħUuVw�3��HA)�,QK ��Ʌ���G��-�y�9K	��x�RU!x铌b7�倐���2���`����w�m�3킺ݭT�dS��m�w5�)�U{d	lgǐ��)�� z��۔���Y�m\}�g8C;�[�c���֕
J��>v;}��u�c�9]���"�E��'j��2�#�ꐀ���3?1�m�Z[,K�f�;�7f!.��dl��5Ol�f�<!q���.��Zӊ��3#/p�ݹ�i�l[��
_̆��1;T
x�jV�a��T8���Tٖ�TO�-馥�����]%xN��Sx)E�X��&z�ݮ�1$M�;g��(�Zow6x�A�Ҡ�?�m޼z�9A���Wώ�+(�Kπn��/%���)>��B]���)�I�,��م��5�^�O3�2_����<�M�؆r�5<D)�Δ��:���J��2�HΣ7�||��2������ms��"�a��Li�9z�r�j"L��I��D�AL7Uּ9�$CSЖ_Sō����u���P�UI�!/:~Ui�%;RC���Ϩ�m���c�$��n�U�S�X:�����1��VR�ȕф|�܅V�-?��	�>�.�őv����� ��r��~�c骶O�]��?sn��~�).�j�]=�a@h@P��mJG����7�K9�p�� ���ھ����E�*��!	\��%�-`��;�u�|�nW�+b�ĥ_�*� �#�ć��T;?:�l�Å��s0y�Xy�b��X	s�I��<6û&,5���
M_�e�����r��Y,�E5K�s�wά���ڃΥ�k���ə
�-�1
S5���&8�N�<��9��f,f8� �b �j��s?�{���L�P��z} Pm E����ltlu����n/���❒ߚ�"��ݱB��$��]�B����U�B�#����,G��C�|��z�}E�k���95�E�d�"]g|�#����}����g+�r�'}�ڠ�%e%���[ą�롲�z��yw�L�!6G停P�-b} -�}�:u��1삝p���=�$
i�հʓ�ƅ�}�s�PeA(�w<�,<�����{kN��֪��e�'�[a��xוQ���j�N�#��^���C*� �%�&��C9����)���EM:�k�/-��U���^_���Υr���'N��8�G�I�r������`���.��o(<Q
�H4�^ɭ��KԞ�A����ߡ���?����0ׁH��
���7�=����/�޷�m�8tf��v^<$X���"����Ct.�,�g�շ@�e�[Sv��LI�J&\�윤�k�ȸ���fc�x|jYS����h� �+�X�w6�Dh[H�d�+�|�|8�/݃���O�8�vS|��]�"�$K| ~<*�jz��to���"���(�:"V��g�7a�!(ٱʂ��	Ѕ�I'�K3��}|��g�S�J��(�Z�أ�\%�T-W)�Jh�٦�g�ІJ�()WxL�G�b���j��W����o�w�!w*Nγ�bbo7� 	������i����qn�aQA�1Y5��rPV��#��R�"���F$њѫ�\=�%n+v}�c�]m����uV}�����r��ǣ��Q>$f7�ȓB��g^0�[��M�V^�4f_�pdtJ�i�NX�C�sE}Ă�6�ٳS삹���H�̜�o����g������9I};�����F�;�?ֱQ{��N� �#姬�����AE��p���M����K4�"��R���|�9i�=��ʋ"�T�����K����{�W��(r�� ��+�xh0`��Q�*ٜ�=�4�yUs��<D� ƽf�>��>�A����������6��e$�4s!̅&M�v����ҵ�R��P��4-�y@;^�p�}�+�v�4��7N��Lø\0��H��i�{=T� �,ر������ݩ)�c����&_ס���3�v�MŉF�i���e��}�w\��:�=��v�}����
1y=��F*�A}0�Y�d.]5�/����0�ݞ��y��A�4�@5�Iz'��,�G `f�C������4��>S،�\���0Q��3�w�*�A��)V3eODs�����
�P��s�i���pW%y�渂 ���*�,p4����Ht�6�m6����W�������ԅE�C�e-�z4���ə7S/�ڈBV�Q��_�r�zi�r�@����GG~/�H������{��;\�n��~BhW�%<�K���y��s���k��y�%��i"�W���.��)�QZnkO�@⻄�F���l��P��f�8�j�n�-�ةDI�ͼK6�'���2��~�V�?[�8�5�ur<'��R����v)��I�0r�� �
���
�?c�3F�H�/�ɽl��z=	��.�$� �������9j�A^`���ޢjK��[�O+���Gg;�N�0��pb�25�����'���P��1l���V��ϲ�]5mɋ&&>f��h|}��C�m��5�0��#�jR/�ĦB�Le0�;D��ÿUỡ��aa�(��Ã2�-O�e���=ޒ�/w_n�T�2�i�~���9�$�k�gg�����V�NƠF*�6�̢7����2S*��|u����ϓit����w�7�O�=����d�;(��if�>���)����'�=���u-�VJ����ĚO��)4=�v�h_>��A�S�kny|z��M\�{E�������1�ґ�PS�_f����6�� ��\�@<��B͍�u�������=�{�T�s����U8>�C�F�{a���Q�4����5��=��+U=��6��onxޝlB����oE�웏s'<�X3�;�Ē秹��T�5��{[̜����=�	I�Y���B��H�����F� �B�����������U�8��w���8D�!�)ˌ���������TL@���0N�Z< D�߆oj� -��� ���ѱ�����~Fa 4?:�8����5��J����g��s���J?K�Ŀ��İ�`g�Sb2��b2ߖn|�]��e���]X�DG�CtY�m��[����&A���!��d��lks��	��:�9�%�ua�y��5����>0��#�	���Jia��28�]R#^���-���j���P��.��&�F!H�8S��n!��2�a.�5Z�|6k����/����z�Z��ⰹ'��H
������{I���RGС��Ҙ�z}��,�;���rg-��-c@Nqzo#�l���	=P��?a���N�Q�w���͙�2p[ߢ����gu�l'�_�����yPc#��x 2�"���AB�P䂯`b.@=��b!�#^�r��y��Uv2���ύ]�)�-7�ÌՄE�����7�4����C�k[�c�>���!%��Q����~X����F�w1�㛷�R7��#�(s]��2�_���x ����H�3!.#n]� k`���.j?�B)���BL��Q�Y"��[1�{볗��D�,�f"���s]%W�N#���>oЋ�e�>*��+P>+���	����wy�/�(eK�[2�����$�����QK��=\�f)��7��p�^S��mc{G�p��8�������c��(�A y7��pxK\cpr
:���6�{O�k؟Q1#wd�woO�o(o��I���������������8WW�M�i3o������7I|�F����X��4�@UB7�����R���[�ԑx��Qk��G�Қ\�x���2� [�k�]d&��v���Km��5c������=ӌ�N�VL+�'�Ý:��!,x 8!��( l��Q���k=�����k�K���O�녻E��8[�%#��������~����\�E��{el���l*} �|R�%���\zo3nq�$4;"��5�	$����_��jk�JG���H	� u�¬�<��b[ښ1=��Ip�,	>5�����J�'���۫Q���ת:(��J ՛ʚ��P�0P���B6�_I��(?�>3v���њ-�}�J��MF�L�q��~Ӱ�Jl�[���sYz�$�u��zJ��4Y�h�Ȋm��@����@����r��^�}������'�C��ނK�)�k<����zj�0a��_�����/��>^9�aX?����1Ŀ-�=^�R��y�Ss��/�Q�Tw0�}L�\"?�W��������1y� �ğ�>�:Q=�h"�:�	 ��B��C��{p�����M�����M��4� ?C���M���]W�&�,ǭ�vh���N��P�����"����n9��v�����]��~���	�Y��7���K��r���h���)��'�.NNm���a����n�
�w M�U�S&ȱP�j� M2wk�sL�3F4_��1��0�����c3Elנ�s��:G_2�G���ö��[�2����(���z�o�:wic	�2�mmM#�[?S#���^��Я
Ê�)b?Uw?�0F���Sh���*��[܌k"$6�������K�Ѧ]�Pfr{��}����Kv���w�� B��"I��3.z4}�gs2���'�v>$@�"�>�˃��D;��;��jT��#s�����Y�?��?�Mz���$ 1�~/`Q�v z[����́�S)����[E\ݹH(ֺ����r�e޶<��2�j��axXp>�S�8�Iܙ���ܷ$��e�ke�
��CjL,݃�\+� �ϻ��ی���(���d7@�܌�s��2K�N���-& ���v����;?2C��\��70G����NX,�ʫ[��Wg�[u��:��2��x[�s����F`���ʬ:����ֈ�F3�	�c)=s���e���+�f�_Y�����Re��)�Eg ��h�'�5���w~.�#%n�D�J���U/Zj:/�&�"��6�i�!�!O.�;(���;�ͯ��vM��i�����5	��E�+[�5> j��9��w�拊V؝]��;��ű5Y�
��'u�����@��"�'�Vܤ-WV��F��zQi����[ZQ*di�C|� q@�D����$0�1�'qߝ)����<&.->�4�e�o�Ӌ���wI��f�¾c��ڻ��c�X�ek_8&K7�O�B��G���|"��G�E\��b�axd"?�A�Z�%UwTGiI@�2��޷�ߢ���b5���G.�FD��W�&Y�n�_]����ۡ�֠iJ�8}=�Qho�^5 Kk�}agΘ��ܼm]��VS�����G��������}_^.������������P�]�|���0G�F\�(�Pe@Zh'�=�/�v�� $C� �ny{�8���9�a��jǤ�y|��EW�.���q��o/;EC���[P|�M[:r֍rV�9�v�<�yr`��X��%�r�`",[�G���`u<�������e*,�,V!x�>�t[�Ji���q��*�b�����7;چ�ն;���V���r�7ń�׉�T�)�a�����9�#�Vۍi�7�*�1M���-�K��N�'o�>�9���� �[��~rI��B����Z������S�z�%?qt���
foF��d	��ػ��n|;�bw�ɹ��3�̠I~��i�7F
4�p��w�����d��h��(ɮX0��#�Uq_�#�6���p~�D��W���)>n`77��j����ҿ���[�ӕ�&����Ő�"-qzn��[�,��i��9�� ]cM��v�g�
��/+}~Y�K_��$��D,���?���>�'�
�3K�1O��0T�"��\��e�O/��z�?�����V�d����c5Ր7�0��Mw@�s���u��x��O�d'z/�'�0F�~Y�������t+���~	]���dP�����}�0y�uN�_<h�N�7s�|��vKe!b�[�a�A�7)%�GXiV�$���v���.&%𔁚�Z*��>;]����.�2�#�z�rrDNL�bJǎ�{F2�Ao#��Z��S[���f/��<���~1$�Y77�b�P�p��U ��}m��n2^JqS�6���v?�8���1�L��[�=�����%�{�Y�����S@�`����,ӏ�cP���h��>�ɢ{^���q���G¾�L���/H#�D��q�QP�� �~��6K�|�P�m�}�|vٸ$w[�ʓ`{q���f@c�<��YqS�7�$�����[���a�.�S�~�Gz
��Л��i��ܞ���&O�Ȭjo��*C?UI�):, ��n��y|�^�����n������,��6���K�@+�wN��?����y߮ J����ʍ��&�l��O�Y�^<���)р��_�o(i��|o�WEz�~V����d�ef9l�|w�4J����8%���b]?f��,�� �P�J�/v{���Kk�LW�f�������[QG%?�X�H��1��6b��y�6���r�%",�ᨅv7i?FZW�+����Fb��A��D�zc�\ё�a_T�!��D�`jg`t$� �|�>�.+Ǥ%��S�9���^ܓg4�e����Ur��]��kxl>xݹ񥍾{�>��AE��i�:S~�.�^�}q��v(}����i��c/�_~��}��Ó�klۘ��Ւf��mP��Gs�[�#5���C����������L�����A�S���������<uv��x}���V ����e}�g,a�-&U(�wH�-�;���?��^�%	�/����A�Dؑ���-�)g���a0�o����Ǝ����`��\�x�I���c�/,;���`���0|�X]��E0o�� ̺a�y��N����2x��/Q�pN�ѡ��~A���a�-@�ZΘ�MΗ;(?�#h��Q�93�s�P�Ke���<j���Zğ��W�ӷﺡ���T�Y6�4��Q��nΩ"e����9�&��GˆC�:H�f|U����Htny+ӳ{o�p���+����*NG��\�֓�	���Q�1h��:��Jc֛،���VQ,��Z�	�-R�$����o`���m��C]-�hLSCR�g��c��`�O�d�y������;9iQ��xS@|o��k3;ȓ*�m�ʒ�����^-�[����L�<�Y9N=�*�N���4/�Ѫ����G��S�d��z��v���QMo���Ҿȥ}~�冠kS³�7�|�A��cê�NVJ��߂���Og�@J�N�\����X�p��䁆`%1i� d���zx�Ήz����e�$wӥ+����_����k�����v͍?Q#��P�����d�@ů{=9XX��|�	��5^�-�������6��^@w"/��g~Jq�;�y&82� �v�%4���w0j>߄O�E�+o����9L�?��g�N�p	\V��yV���)?������������W���i�-� ����EM�e�c��G�kb���J�Zt�N���z��U����x�')�y���z�mik7���H��p��#��'Y�7c�3��l#��J�G�HDH掗�7t��$f����6�(
S
�A�=����@B�^h]��T�^�B����F�f��ج��j�9v�(��> s?<���Z�yc��g�g]�Q�W���s��ԏK1�N��T^�*O��'�^�snR�v�����@<+�\
LE���Nަ�~[?|�c}�D-�]1/}0�0�M�0RR�1�$�m����2�£k%?�������iS~�Lt�n�"���dj��3?����^��~4j���Trz�$C�pre�Gr��矰�{"a��Z���{�g4,�ꯔ����ZK���Հ���/�G�Ez��P���M�-�iz�o�����O����"ذ���τ�x���% z�k,���b�&���M�6����ej�d/�[BR��K��p#|�@+��*y邳rA���|��٦���>v@M���S���L���Չ���b�@��v�K�~P��m�8�V2����[IWڛ�^�������JaA��UU�pW,�߉�=H�V��7
�+�_e�hx��Ws���(0���Y���US��]�d���G�[m$�	�\�
��Ew�q����ja��V���ؔV`��QA�M���ڭ3ׯ�s?���P���u�q�e5��N���";��k'�mN���r��ȨGWS`� ��Lj�.���=W��ǁW�)|�$ߪ� �&�X��%W��d$�9\J��CP>��~� �ֳ��[�X�˚Ð[�����7?PXet_&�b|��p��z���?�t�k���r����s6�M��(%�T��w���Vjο�V�J�	�b&�B�Eu�u3�J7�i��D"3�;/Sr[��������=ZwS1K��?��'��
!�<l�~��d��|��l���>WjUc��eg��1�� l���a�.R�r�y��8���Do�C�����]�º����O�pV�6��~�����x�y��}�R�e�L�=}�:W�G�A���+�m\ ���9,6�Ku}����5h��QM&�R._����Fߟ��)��xj�Z�e+Q�3�a��D3��a�f�?QN�Pi*E�9��4������Z���H�ĺr����<-���(��?D��ӳ
#�\?���yA/��i8v��v�S�CW`R)��J߹�xͳ�����FKs����2 ?��� �{��b�3b(�v��'��]�!�2✴ȍj�O�`��"�g�^����Z�l�&��gyA2��|k6�Q@������@��	��a�rO��8���MF9�L�G2 [��98�瘇5#���i�=��T�ίT�E�\�؂���e����ߪ���6D�Juyԃ	�eƏ��֯�Ϻ+�D˙/4�>,c�\3��r�zd���M9��!	���S��Z����>����5���\�Z؉�n�w,�����H�s�3��|bZ�B�3:	_th$�?Su�y$�C@��#�*07. [��4�ReԾ6���w���*�� lQI�~Hg��t
y@��#Br�#���Ay��mp���l��RNi���wJc�'�ؚHCV��NB�MA} ��=|K&�qã��۷X�(�ƫ\����c�?fZT��T�?�J�l2�p7`y����tך��P�M�G8�^,�K5���n'�{s�輷�T�W�������Y�7��Xc1=��n��E��Ԭ�q��H�Y�9�%Q{D7�F�!|��>�����k1���s�g�ܵa�fdcN�Q.���RJP^���22������
��t���S�HW8�5(��?"{(<{d��\�>�Z���"�Ѹå�N,�6��\���UP���%�w^���?M/��i�r ��%W�p�(h�_}�|ɉi�k�3�ww,�[I�2����E��X2��j{�4x���@�j����)@&��O���;?T?��-�ۏk��.4Z�CN����b����5��X���l�*�����uz�bJLvr�e�N���kS����w���7��!�0�]��ȬE�Q�]}F�e��	:?�]2Ea�,�+������Ո?y��\��Ij�mr�f�nt\��٣�"�;�4[,���QZ�Xc��o<k�S��+�����)N^J��>+y�#�t����� �>��C%&@�W�7���m�чm��������c���Ú��*���;u�|@����o�kT�^1�01����fE(�.RBT�?�;�6��3Ɓ��s�H�"&��F�ubh�E�s�@��1��X�כ٩imh�]�2�"�Tl��#[+����R�#�1f�FS�~$�8ty�qF\�0f�텎3B-���d����H��x$�'��x\�[9�b���,�+��\M�#�ۘ+�_î���/+��f��"��EK�L�B�F��E�j�t"_�$ͣ��_۵���>��u:��7��J6#օa{�N�z�[�ƪ_���hM�`�NIRE���u��f|(OBW�9g��Mj���0xO�x���,��=�d�J�A~5�����e��J큦E����D�Uk62�d��N[=d���C�}�0�	���r�|#mذ�����.W�}a9��Z��u��ae\A�y{L����YɁ/�&�ç8�/�C�3Lt�%fCgՉ�������`.6!m;MT�L�1Һ~�z�~�>�&�vY��1{Hi����n8M-�!�e�
�uQ*v��W�8�/o(@��G'X��* ����wD�V���<���tE���Z��PM���V�K�G��Q:ȎT�7v.�:ߒ����Y!��*^j��8�J�\f��0���ߚn�
V�W*/����|s�ŏ��"�sPK�z�����&E� "��p�嗴7䋂z�4���p%ğ��hص}�0�a�#*6,�_�����@�A�t�۝�є�OMdJ��V:�>��߸yH�=8��0ǡ.H��O��"c$渦�>�s>j(T#>�ё�;c���-��=�[��uѽ�F����_�|Io����yo���|����4��7���l�5�] ����V��?�ö=ŐS:w`�a ��>����g7�Q���w���2��R������U�ݽ'B0�#9�C1�n�����\s�2���s@<��
�P�������jD�j��#��#!���QF�����T	�~�t�<"�o{\��K���	(�aW/6:��<Bd��b�lźh�ŏښ,�Pb5�v�;��'�<�2�߱X *��`��;᎗-V�ƒ=�s����&��=Gw�����d��,�T� �\�͂�ڨ���Lsᙝ�AK��LJA����.����^U`��*1>�9�J�f��nh6 �����Bs{�;j�����h�%{w�M��tl<�����u��� b4�Oǰ(����5P�T��lh�%~k��*�=��j(���~H(�sY]�A�
��8<d�t%�>����VP�̷�9�8ҽ�II�I�i��mh�{r7a��H��&K�p@ma�b~d�⮫�f��eVḍ}��a�[?L|
��zZ�����s��{E;6�b/e��x��%!+o�$i��[�����v���ɓ�4;���A@i/Pzw=��C����S��<q/6�B��k]0��RH��W1�����R����Q���k:�d�F;�|�pNK� $�����.�b F��\aCP\�oM'���ud����C��-n��U�  �$�(����_�5�Y~��`K��	��t`;SCB׶�S!���?�JHk;�aY�X�89��ʐ�V��_���I�E���[�;�:L�K
����Y� ��YcL��:^�Rt�ײQ\�x�SKB�	�]�cTi�/ZN8{8�e؋2r�5!�Jw��3b�y$�4Pi�l0��@�-*r��-�Ƃ}̹���B7�����T =}�+86�a���i�6U��DL%�$V���ǣ�����5Ι{%�+H�� ��������#�N�9����&�����ࢨ,�:PL�v����\$M���dҲ!(:u�l���7� �w"3=N�Z�noB؛��1L{�)C� �����)����o�Z�\*/Ϝ�j͓��wY�}=��7�>-��2Ԉ3lm穉r��*�r��;��,xFE?�=��@�-�����v�,&}!���%�����KO����5[�[*���b/Ȭ����H�G�gT>��U��4�H �U�5W���?�Q�2��N��	�w(*��f�#XZ�u햝)����2�K,�jF��J�*��^��t�N@�9��,+-�g���P]Wh�i�P�n����6cFly��'��ڐ-0mȸ�Q�": (k���f�i�F��UU��d|�"B�6�]U'&�&�0�WM[�d~K1�	����X��~h`� �����
7���=T�<'���9�p�5�Ko����o褪q��v��@S�7qCq�=+��W��֚�D��aOX�ٲ
E4�P��k�3��� m��s(U�]�x��1/r1o�!6pūA=��~k}ǣ.Z��%��wnuW��{�'�����Nݻ8�s��!�mꩾ7�#.��4	H�B��@/����e�Y��L�")���q��;\�K���Eߣ��֟�tv��.�y6����ͱJ���oq��`�j�k$ŷ���-�p8F]����J�33�������-gJ�rM)�_�	�p��������C��[ ��u�*��M������"�M����{g�$ˎ�N�>���c�dħ�RĒ�1�;��+���_�\C���Ɉe�o�!�T�.��G�<e���p����8��(J�3t���A�S�����|P�����%�TPU!�S(����خۧ��6/���N��"�L�s�,�B�Z7k��J(�H��o���_���r5�.N���I�������r�V'���7)��Q�o�'�p�(����9SHSǓݺ6\�,-w�=����JAqm���E���H\�{���Ӳge�YB�芚�h�e��l�v���E�s����_`�:�S�����s0�d�����?c�u�ኵN���WK F�{	�"�jga0�D�œ���)�rʀ�QK��V��\��d6���ő�}vU�Dx �Q�dTBԲҗ�5ֻ(��#a"��,���ʘ��J�8S�Ԟny��$<2:�_����t�� :䊆��f��!3.�	�ߎ���E\MR�ٿe��v

���j�U���&�[��Pi�S�0��@���J�zq��9e��<$~�^J֫ό�s�q�yV��,���Of�8����W��	�D��KH��� ���!2D�[K�4sJAV19oUT���ۄlB}T���h]NtB��*NH��%#���#64{��P���pY����~�nyQ�f\�W/|��v�/dy�n=�ң����s�[�}�`^2���⟫b=/�vni Ĭ��Y2N��4	XI����-�'��p�%���Ǿ΢_�TZQ0��۟����>�o�fh���9R~�>LW��:� dz�ӯ2N��!b>I��3��m�-�D\�_"!J-d)X��@kd�G�M�w*���ws,���;]�}5GƕT��	v�%P���KB�M4����6;qȬ4���Z���u���g�t��7Cƞ�y�&�闃N�R���P�jL��d�wd\wQ��Q\侅}*�6��$�����5��꾲�+g���A��c���j���͡%m��M�jY*�0ջ�}�)�G��[.p��CHQJ��W_�|M��GS�h�L�����h8X�����@V�S���B�Zݲ�>����͋!��I��ʋ��q�,,�c7�A�L5\��CHIZt �'� �w��R)�)-G,nۈh�����f�~o��K����<�#0(+_
�X�֗��*�H���`�d��h~�e���U�Z��%�#^~�W{ʆ�o#�
X4s�,�c��8�l��O|Y,B�J�`A@�}΀�	=K��ײY��K�<�dާ������
vC��#��[O��BRw�^���0͂!��q,��q�H�8�� fL{��wr҉#�ͽ�C x�޹��Ϲ�TJ���� ���uV��+O�  �F�*#JU���e3������g����o���GZ�������=$E��Cx�:�3w?��iH�nN�U���'dH�$oޗr�P�9�ǿ��ns�'�M^��A>oq��+��{L�Aę�!��i�/��y�ቾ��p����H^x:�����L�����(	�妏�G�~����t�î5�e�f�D1�$�|���u�<ĞTǋ5�����#3��Bюk&����Ͽ�k�zU��5��.��Pˌ"�,CN��ل{Һ�/,Kjk����g�O�4>��\S��|~��'*KyY��:���CDm���+�[�߮��,����b�ŭS��<�ާ����Gg͘JM���o-��B�Ġm{��\vL�������J�L�2>*:�L�@�d͟vuv0 ��mP��9��0�:�u��!���Q�i"�گ������YB����� ~O����a,:I�!��M��$��ݛmz�Q=�gKK��J�0�K��#��f,�����E3Bc�A1.� H�K���%�'.{�ғ�}R��@ģEOb�R���MǑ�d1K��qc���m��-��nk,��sn�1@�Mi[zX#ޒd����q�y��cqP�6��H�۸�S��`?5b)L�c7e-y�ֺP��0|E2���H���OI&ԟ���y֧�o2�����~J��5I�	�"�q��˫Z�D��FPa�q�p3���4赧��9�)�QN�ӱ��l
���%ө��*-�j����N},�|�<L��t2�1�1�iC4`���G{��\�'����e�����E�Χ�!�V��o��@d�K����	P
n�M��v�љ���r�+��^���:� O3����((8�]�1ze����W�Y���#@\|<�9�����Bv�$�� ���p�"�Smx]�a�����Y�`hH�|����'^*���Z�i��񭬝�ZΪg����_�;��%|���.[?�X�f�*�%��up�Ѣ��\�:5���e'T<M(ɭ���L_�pUM�n�x� �Ϥ�z��~�%!�^���϶��)oi���
��tN�@,� v�*�� �&*Oh������Tr�-�m�qъ�L��ZC�����M���uͿ�����r� 8�1�h�y�+�O�oYu`:����㸕0��6c�W����_�+��|Q�\k����J�����z�^�d�-�'*�,o�bM�������b���А:�7v�ఈ5�+���w��_�6��(��e�½`!1�c��o�hh���+%�)1֥�bW#�Q�f:D�]�>(��̦5��
$�ׂR)��[G,.�$������ٜ����O��g��C�+P �����q��YR
|>��Q��z�m1Q�Q�����������p�E��9I��o�B�{��~�Y�O��{9d�VKd�k<�%k�6�ZY����-v�$��OP����2L0�,�a�k��Z��r�.��ocڏ>��Tj0���+����A`������|���_Z���e7dpG��,�Կ�7�Uߢ�W�Wn�_O�{,�`��}0������ �>���:�d�o�ʬ�cs��2.R3�>��Ԃl(q����/F"Y��1p�`��� �s_	n��2Z����z�����_D��1�h�9�1"_��]�����߹� Ԙ��W�t��\��P�ړ_�R�	ì�5�Z��b#b�"z�A|��F�1�#eA� C6��/�w L�Ʒ�E�q��J��Z%�R{� �v'���A`?��TsZ�>t3�2d~��l��� Yg��@n����$l�*G����Y��<�x���!$��nY���N���~N�o�K{jƦ��N� ��yQ�\����z5 :;��j [�7�u'V�j`�H���*�]˂��YB����z�f:<�gv�O��Nt�D19��k���׽�S�B���d�!�3@� H��p�}c��u&���O�=EJ�TJ��(��٬����)I��4����h	��{:��Io#(F�.I"1���H��Fxԉ��'w\{c���-��J������)��>�ZC2E9��@c#;�n�.��d�萜��,�js�t@V�͓�N8����<���z7��:�!����]������ϙe�Xgi%VI
�� P�Gcv��[�LU�?%E���S,�l_�E��|S�<��1���78��-(�N�8}�ʻ�j2+�Hv��D��гC���쏵�z<>������g�jQ!���o�V�o�����>����j�U|dvR^ʜ�mAˋ�l�����8���&L�._*M��B^f��Z�Gj�s�.[=*@m�#F�}c���
��� ^�ZM���.�a� �	$�Xb�梶	���z��W�:�t��Y�@T_��|��6��HR���^�&rwbo��G�AJ�2U�+�J�{��F���Y�a�!��S�a l�Ϡ�����`!*?X��58yytkhkz�?}ឤn���5]��D�W!�/r6��M��$um�R�iLĖ�X�L,�y���{��U��wU?�A+�7�/�H$�AXqj�	[x�9�n����E�dY/	/&M�%jܜ�堚NZ{�y;��n�`�l[%�)�E�z3	1�5\���Cfk��m$j9�χ�,;�1&~�x��b��l��rZ>�$ED��ޠn�Jwxh��]Z���`��_�r.��Z��b��X����,��Qn3���ʛd����1-������|96��ge,����ZqOG)B�����lT��S[��A4W�K!����δ��Ȕ	O�n= �~u�ȩN��z�V��&2'Ǆm<�����DoZ�h�������-�W�s���IBl�4۾�?e��soy���/N^�@���0�Ք���s�Q���Z� \Ǻ#�𑦡Yٓ[�pK�O,Z��!��H�1��� 4 ��o�9˾�L.�����%{b�(���ɳ�B,�����Ĳp������8!Fq�d����BBjTژ8�dn�!��)(��sgoo�J���q���p��2�BY��7+����E[@CR��g(r�����.���:�u�@��T��KPR�.0�z(7����#����7����o���Jf�.3ga����d�������>$����-�*� ��=�����g���=�	/�u����{�i5��3�2����A���q{��5�b2��U+��1�ޡP�R�͞��%c�ޑk��КY��U�ר�ؾ�5R�tm��)L��=�ea��(��sc9��},��G�Xb��cjx�T��%�~V~�v��ո�O=-�v�v��u��l,Ѐ�@��%������#�b83n���7��l��X5�2n�[��u�>~��r�;<�}�:{K�����=��I��6��Z��[�T�e&�C��iHh6�n�P%����i2��r�U� 5Ŧ�N�����u�˃H�~�|,fU�	�!��|�a�\����v�5�R��*m����JH�Ul����:4��b`���3z��l�I]8܌�n��a�xZ�ѷL�r��Z���^�j�h[�:g�!��9ʋ���cC1t�p�����c�'J$�U2�߹��n$l�>�-(��T~�����kq��B&���xpɀ�'<f�ʍ���S.�d��J��0��)u��﮽��E�T��3f�?#�H���u"B"ZxY�7�dm:��I:�z;�'��6��Df	������y=�ʽK��2���d���%���iU�
R��U3��k�������� ���^��'ⷦ��*��������s�:�9f"�+J��� ����z F6��D�����(�:2���>0,Xj@`�'��oN�����hV�����d�4�����a��>�:w���}֣d����x��s�1���<Y�N���q�<Y/g��������k�� Հ�*+�a���lU��3	�E��gn��"TW��ċ�P�/%�����/S�����#�Cc6�Q�� �`\9�m�c�&�Mj->4��Q9��w�y)	��r�R&�n��<�b%���H�	J�޿�>"��8'�
{�TH��ܦ}�bQ|���c�wl�n�kj��6v�Ֆ|�8�`��8��,ɼ5�E�iV$c����~�v��8��u�@b�=��/u�A&!�3�C����L��Y�6b[.��r�;��*C��V����w"��ү�������hl���ը�fB�g)��,+bG�cؤܸ^I��ːх:���NsS'��q7Q����uNB���o���<@�����-�m[5x���,���碨�(�zZn���p���[��FCf�C�b�_)��A�?ϮXaR�)�s�ӱ?x�gPK�TRc�,��E��g[p����#�Q��C5e�Ҋ���ձ�j '�=A9,1}]�l�.���ӟJ�L�$2�PϼmpR��=+SF��N��'˂)�gFC�����Z]ʁ�p�߁t_7��%g�����Bh+��sK5�}*F�fHꕈ>�-!���q�5q���<=_^�-��<h@Aԋ�=��8�G��b���5/T��XwC�? �?�������Y���/�=Nxg0�Ҿ�ӈi�r_��a�l����t9��hA'��JXuB�޺���>� n�O1����d=,(������e��g�l�{�Cc	n�ID{�[z���7w����$b��}?3DgŢ�Y�c߆ז͏�84�D�Ee�D�P�&~Cե�c�)����¡���!�� ���;guF�i٧i�j���`��-�^/�9{�NFVC��ַN��P�]8��vV/K�����=�����"�T�\��R���T��̀\|�"���l�e�<�k�.0�����.��7+'r��ax+닡1��H��0[}J��@�r����/�����=ӟ䖏�^+"�S���3K�XL�t�>�YB*K��"-��L�Ku�;�)��V�G�֦)ȟ1�I�q���~ǐ�Z�����H!е���-v_�d.z|#�A���Fͮ��^s���2������\`x�j2������W� ������b��Xs�*" �Y2�`�������a��șd�4��m��Db�����)I��Qwc�h�҆?�6Y�{�������%�/�y�k��E��/�v�ޱ_B~���=�Q�
X��Z�*���bݨ�T�D���<vP����nW}�t�X�?�0$e?<O�)�� |�-Ʊ���1ʏiؼ�u`�C8zߍ�W����ʃ��2o̡��i���.�q�z�c������?g��-m,�\���W:��6{��y�uR{esI�0�ci�l�����GF��,ԷS�!v^�ӌ��������`PJA�|��W��[L�66��0X����Ev����~������%��%%�G�.��j䵏^6�g!�o\��Jd�u^���&�d�������������0��
�Zl�h�)>���[�,�󾩛���wdy��@@�,#y^�h�nwg1��o������Q-!Ze�|}��������I-��D��w��!��wTOH,;}y���g���_��jE�1,G�d���7�Kjv�S�]]��1s�޳��E�`@,����&�{N06a=`������V����`��փ�ш�גM���ʢāqN�>�V�I�t�?�5����(م�K0�����Tr^��<�Ё2�;*P�7z�~<��e<G��A��*��10�%AFJ!l%��o���n�u���$2⾾�+��3)�m2(�n�����Z�QKԣ�7�8L��RH��NY��2�<�:��Ӝ�2�BÜ)C�� ��PM@��=Msd'���/D�Y!�+�l_W����Y�gM���#�EA�D�f��-üg��[�,g��k�W�o��#���W�J�)���"|�&��5r�)��$�CV��c��ENy�
쨨^��?�D`N��}jew�&]�l�M�c��&g�2(�&���Uz�C.W�N����^�[��y�9	w�L�Ǫ��BG�8bxۄ���)�����'��ć�
��lИ���3wW���}�2���;.ϛ���*���ךo�k0��4#`�8�S&F�{���~% ���y߱�ߎ+�\�%^�|]x`��=e7����~7*g���e;[^N�G;O�NݧŘ*{q.xz`�@�z�~�t�;��e�;�P�*� 2����0��<N�7�k	�u>��#�8ݶD���Ӻu�����AG��!�U���,�W*A�|�
!���:�z�ӗ0�_)Ю�����<��3>
�	��jB�'b�*ϴ�Z4/�Q��F�P"�z����?j���=��H������v��S���[�O��}Kw��f�0�I
�#S7�4�2`�d�!r�`�L��[���VK�2x�`��8�H�4F���=��m�'�/�7�g�n�H��H%�nt`���,������:��Ju��!ߏ;[�|w���.���Z����O���+<:B���O�B������]�ٗ�8�|����3ouI���=׸�i��E���&Bb��$��Ԫ�(C�߇�ʐn�
%	�Nw��a���j�i�������y���d�_���d�>�"��9�Խ�(��WB�nt�=Aʈ��-�+�q���}:m�#
x��SCm �ۑ���b0��MA.;�P�E�~�m6����'���u���K%�-dbZ"����c;p���6e~ڽ=�����u`��kʺ���re�2e���	��w��l�Ff��`F7R�6#�$�y^�G�!Bڱ��h����Qv�9夎߲�qcS$��k�
����&��w��P�Ȧ�pJi2��'�P�"0W�{M%�YQ�]�B��x�����W,�aK]�%���#�}F��Z�٥t|�]��t����4i��5`S���_w�|��^j5�9	9\oevf�'�z�Z�l�-c_w��@����D>Xd4���\>CI�c�@�M��G����P���N7:O�o���"�&�j\�">��1/���z���ȫ�>�e�3L���N,�GH�������l�Pμ��e甠�@�����#��.��THN�d���9���v�|5Y���}��a�X�f��e�{���IbK	�K�Ԍ�~K���ħ� im
=D&`��~�����������*%S8j���u�� �I�6�D
��^�PK9����M3w኎*(U�'����tU���r,O�[`Ea:�|��%w'M4�K<��k����_�t��m���+��{Z�����?�����85?�~<�PT-Lbs<�b ��gzڢM`_��?3Uv�X��?�7@����'�p�w^�ǄD���-�W�e!Գ낫�e-�5q�g{i�N�嶱��R���+�|N�$��|-%��6'��u���}�p�u���K���RtOP��y<���lt�6��{'�˷��G�~�fr�`e!�Xۀ_>dDHI�|�O|�v�ŗ6�)�� 几�����-4͑Z��/��,�̑�!��t����4l�C��X$-���Pw55Hfb�Aq2+@;u>��T�T�:$Lp��3���㈔���Sh)�:&�[4ξ�FY�y@I��'E�V��{���WQ�SYc�"��@eZt��n��TiŘ2�\P���@��X{�\��킒�EԨf� ����j���[M�R, �l��-�)�3��[h&D}��;,N�s���˥���sL|��hS�8�W{4K{ŀ�-h�@�yYO9�-���Lb]��[���] &���E-s�[4�厯��8������ZRi*V��-� ��/��_t�9�����5Z��ų�����,��<K}Ӛ~:i#w����`���d�߲��1e��k��2�y���4�����J����'	��f��'���|�N���m��#?S���z�����OM� 0�����+D|��&���#��a��[F��e0��i��wm��6NƱ����Zb"�_t��x���g��V�/0e���BxK��|B��r�^���3_.n**��
� _դU�d�!*��"8I���}K�����c�g��7zz�M{vsS��4I���2��5%{��u:���/�j���푉��?��qtb���doq�}��6�"TE��e���Zrҵ�0ew�`�6'8RѾ�T)e; ~,��S�h�Z�ۼ�2,l��Če1 �:��׌7?��KI%�`�=�[X�oT+�l/�97AK齎t�(,�I=<���&7<2m����?EN
��E�@��6I�p ;"���;�y3��Й�L��u�(q���e�:�,����j���k��E:m�%��o���n�7�d���n=�w~m�1�#>V:��*�.���Z^���-a�r}�S*������Ko����_*G���mĈ�I5�Xkca�zЈ�.���\�jQ���5*��ц���Jzސ��e#���B�$ij�냫�_�ĈR$�S�����q�];�V���$�A��_�ŉ*��i@���EN�t��2<��J0��ୌ	T�db_]F��(�A�":�4��b�٭���_��F��fR�dÖ`���|�Sv�Q�pQ�.��M��nZ�����,vfm�L�� r�t)U(UG����kp>$X%�u��I4׬~ھt�N�#s�����F��n�gN+��HY��:�"�o�b$�r|��L��o��WP��Y/[�|9$��N%�6����0�����~T�	1�o���H�b����L��^�c|/��z��f���#�7��fz��YOn��*��g`�\���*��h��z��k�Qb��x�n~-��{��}�p"�ŀ)�E������I��{՚��� ��_,�r�7�Fn���6G���0)pٿ��k���g8h<y=T�R�{������}^�"���|f����3�| o��A�`o"3zȸ$W���-�SZ��h�L0��
�/4�,��<��Op�7�siџ������H�;�f3��W\�������NNճ �����@�tz�-���u?�C]�=��H���TӺ#��8�#���>����d�b�O�[�z�J��|�ED�q�2�c�v�c�mx�-h��}�x�]:A��mFk����ԑ�H�E�p�Mo������&�H.���
*�1�L8��6V��X:�z�w�n�Kg��ap'��������6�=J[{ւ>��|f�j�f��`�>6�T�VE���$��z�I!�������>�B��-�Qt��3w$,A����r�3��n�E$2V{��sP�`u���r,�Z5�򜹀a���P؉��ר^[���	ɽLg��_��V�p]^�˦�<'���]NJꢚ��.P�p��E,����L��-Q��X֯�<��e}���_;��z>n'_�J}�����)H�#��g�$���N�k� ����3t�o.i6v�bq�ĺY�T!���)m�޽��|\nN�A���6�T@U�������r���s�n�Dr#��YN�f�*������سEܹ�	(�}�}����[� �¬��$�HfL�}��5�<�**�jM\J8q�����PYyF�������4�6"�k����&��,�ı�q�1������f��?ر0�*�u�9�;�N:(�5W'fhr�]�8A����W34�GWR�Y�"�l.1s�oå�P�P5P��������JK��:)E:�2�����jJ�u��+��V#�Qtc�N��m��0��G��!�'��T��(}��;��g�AN?�M\�_���b���jJ�ʃ0q���[.xs!)J�Uz�p�LJ���P0D/�_B;s]Z['�;E�y0W��Ga�4�x��됐Uok|g'ƿ���NE%�>�%9�����K�a���U��PeK1������vz�~�-ݯ�j�GE�joq��rQ�4A%N�U������X�@�"B�k|��bE����c��V�����a�o�#ځ8�v$�c�W����B���QK�eك)exL�PE�ެ/t�ꪦF�g�nv�+"_�I����H��V��E5�t	b3��w��s4�3�iJ�\��ف�"�>}�?����n�MM��<�9F�j/E���
Pz�<J�����s��
n������"b^��s�s�KҠ��§�S��& �B'P<<]&�f��9:!xe�����e�X�R��"@�l�ח�,R�y�{8)��o�I'8���9ٷ��U	#����ɭ���6�I*] I��p�,�B�r���\��3��%������WV�"TNq��IX�v�B���/�\�&ũ��E�b��n���-4���xl�~������D�w�+����_GG�\���"Zݥ�r��٣P��?)h��oFuL����:��3z���6������" �){������.c?������Y4��Ğ/�����,����p��ޙ��(�����PV�w�M^��E!�w���#l[�|w"T���^C�h
�aM��)�n��ҥ<?�&@���9"Px1{ǲ+?*��T�a�Z��8���y(�F'Y���v�o�e�����|

�B�j���d�
7��<����Z�uX{e��Eg�i� #��鬷*��������������\��ĵ456�ޑ�>�Q"����&$o�ٹ
�b��f���Os~LY����P�D�6u���t�-M^k��9!?�~�)�}��z����d;�iy���Fzq4����=?I����G��B2º�"xQa}"�����R�N���:kݨ��&ɲ#�{J
���f���%&-S��������#F�#]:�{�#M�@^eŏ�E�!@��k�r�l��G>�:1�%�5��q'#b�"|��.�1��%͝W��k��7��i���hLv��]f^��kC�b?sW�fn)u��<h5�W�u�EM�{2r�7�����%O���H��j�ճz��aՅ�����%/Q��FG��"��TĤ��6N!���|�#zq. $���9y#���n����"�e�'=�-��2�*H	�[2�}��)R��3�b2a���`�"�.�M܈x7�[��oo��5�/��h�f�1F�rs��T%o2d�F�YWr�#���T�LS�4��DB�~�8K��5I`FA���"z�/�ȩ����-@_�p*�y�ܜ�r�+�R�dٮ�8�s�ϴh7B����V�yg��D�WcqJZ�֭���8�o�:�|�".���x,#mR\�E�6�jsw��������Q���e
�PaU�����5@	���$�5�RE-i(�a(�� yR7,x������AdS�+�Z��sn?"'|r�U�������I�а� �4����h�v� ����@�x^tM�̯�o�e��7���;q�����1��#�b��2Kl��6�~wl�8��]�C������qȴ��֦c�p�~0,�|ƀP���(o�Wܟ#l�%��W�d~Fk�?�:n'�K8q&�F��Ev�}�[y��԰�%��~4m�be�#��:V1�V���tK-�$0d�����\�X]0��}^�������K��mz�Ph�0�C�mg�gd��#��3e�7�lU-�?&���Q��C}?K��ק��i�?GC�z埫::(i5?o�ڵyrY6x
+�%%t�����d�s���c2sEq��a?{��0�v�.�3*����J?���
�޼geN-�w�K�x��Qo�4��2~�� ��:6�@L2O%�j�L�x��dW�>&�����ŝ5���k�����[(���p��ac+���|�@b ����l���X����GK��m(���j��U� �%U�}�?��!M�v�EH�OY��2��X� }b2#.yO���
��{fj9��
(-B���On�YÒ����y�tj��l��u�<��Mo�aJ��5��Ǥ���7`����n h�_ɦ�.tLG
^�A�_/X���	�M�%��)C�1}�;]p.����Zf%���"ı*�*r��Y�8�`���B��fz�m��l=`}Q㧸�ߋ���2K_�(y
&TR�O>ʳ��rwb�g�T �m�C��є��L���B���Ɯ��c���p�hIH���/<�uٽ����5�:M���sS}ĭ��tBo�!�)�tm�� ��6b� ~m�㺸 �)�*9F�#:��c�(B�ؕ����S��/Ix�N@^wA�T)�?底��T�!o>�p���}���%�~ő�|z1���a˦q"�> ��3VM �i�&|l�B��T��S��k�������(=�J�n���f_����WH���$��z���m¸MYV�@TQi�i����]|�]�������0
�ć۸�֗�g������Q���r�=:$%�K��r&ZM?q�h����iY�l�^�$�XlzR�K��=q>$�����7Q��f\�*v2h���=��%�&�~�d
�d�T�_�]���bq2�)z���Y�B:B8Zq��+�;ej1>���<�h�>A�LxU�E��j.4��3x}) ����M���Q�f״�d�hz��K9L���!4��"y��K�.�U�#�Yβ��?c<�A��c�|�gJ��1��(� ����_�\�5���e�!�̠XX��sl߸�߷�o�6�v�10姷Ru��p_ !�[�� 쟘����eC�����w���WU�e�h�����ې?�<�r9��6�P� Kkʎ�d��6�!
R\��A��O%�&o�m�%�,������|�)�?Y�V����#�Y�0H`����ɒ)��Q�CX̤k���, ��5�/�X�Z|�y��k�_9��H]�tY�b��lh
?1��U��>�����-t'(�'��6�A~0�T
+��,8�tD���R_5U�%{T��L,ƭ'22k��0̌�NA�zgS.��['��� �����^�n+Rh�#q�9�4��5���)�-�>ɜ������pY�@�}4�	_�[P.��0WPfz��l1W`�;�q0f�\�.��3�ܾ4�ٚA�c�u	�5s�����o����>�ty�m�R٦t$$��TK�c\_�����W�[�sDD&`�"�b(�3q�q����M��5�$��	�^���Ҡ�_B��XC�����U�.��5T�C҄Tx����O����7�~�l��/O�:..�]�]��ByS�<j���t5���W�u+G<���
��]}�f=�9u��@;�c���-�H�V���jv��jIݦ5���N|���f4Dm�UNN�]�^��=b����<�]r?�y�l��2��6��.)��}-�"/�Kŧ�F����H"^�6ER8���&?23�� *���nqSih��NiwE��ݳ!j�]ݞ��O�n�4v9}�2��]�FHvm�n�r��h�l���Q���UeGWЇ~׋#�$�vFX��Q� �z��K��ď���oN��(o�Sjk&��A��!��j"Z��q�ۄ��a�o 0�'�K���%y�|�m�$�s�ߐ����Q#H.�$j?�ƧFd��	��;r��ƝY������
"cv���>�����>Yh��=Y	\gR�/���b��@��8�u��\��}J�V��խ�l�e�	9�Hl%g�ޏ��V��ԅv�H�i�y�,�`�>��A�n���$�� !%�k'24�z�"5�qvۏI���Zu�Ĝ.5�66흜ОGw���v�S�k9��zn�%�C�`������[�
��rع�xW�<X[q M����S�h���̥�R飔������k�ޤV6�h�*�}��vP�l"�FC7Co	 කwZ���ꋣ�A]R��wqo����C����ղX�JN<��y�X�[�Ag/�7�N�OsL^_�A^`99u)�e��(�2=C�d�@S�v�3�f\����_�b
�ǚA)��m��_<����h?��� ¦5�f�.�U�#;[E���U��-��>Z�"+|�lH��0d�v5��"5�W^������W�a�?�V�&C��{64,�W��lJ�Yo�>^��dȗ�+�1��UE�ҍx�ײ�kΦ/�ۓ�[i����|� �HS��ህ��Uf?oC�4�/�~q��=��)g``����T�&m�֘�4�vg�ubO��@�Q�U�����"�ruuQ�� �7��d�*y�;c��\�Ǧ$L��?���&_� ��<V����8�JJ�i�pE0	Wdʩ4��%p0f'���*r;�:�¾�B@Κ|rՀ��Xؒ�k/y�(�DZ�舢9]h��g�|>� ��R�p��r+~�5�>�(T��:�VtVx9�Z��1�vW�W2_�ɵ�l�G�	+��U�
s`���T� ��~s��:�0���Gy���0�˺F��j���٫��}0c���=Z��������z�ΕA{+	�v��M��Q~���C�LVfu�Iw<d�cD�~e��#�ܗ�N廲���,�^?�rp� a]�k���~��v>�:�p�W�'<�S��vJH�N0aN0�\��:Fb�ӐƆ˴h}�6:��򀴈k$N�=5
����i�9���f�=���"Ŭ�ㅇI#1�f��;��>�T)�L��=L�J'HS��ٴ+�ٰ4S-㓫�=���J����kթ"�(R}3�w16և�J*�zp��J����E�z}�wGG���hX�{���8� q�Jl��v+s���iU⟩\��i�����N7E��A����
�S�)bDAƚ�)	���Mp$&]�vF$r��?���ۓ_3R�ib��^3�����P�������O⚕	�ey< ,-�̴��Np����a��UY�p�~�\�����!e#�ڳ�K�7��!���Q�'�݈1����0����J&�?K�����ZJlwQ�$���j>�hO:���J�k�� ji_䋵.p`Mx����^r�`�%���C�S���'آC
�S�ݍ�A�v�LHM�~�elv�[C��6z�y���"R��=`���2l�d������,[�f��N�QK�.�=y8O�P�ByNA�޶w�\�H����? H:�@d��� �4lR��-��7��^�}������ϸ���e�TQ�Qi��1��I��kf�<̮b�j� � U4�S���kA� �����Z��a$��D�;W�Z���� N�Z�%̜dǿ�NlF��M�>OO�:b���M�O��H�V�[fq�2��ɒG1̈́�ҋ���,t���-x��2�p\
��'=�&��k[�	�WE�Nv�'�_3i#-�|�����@����T�*q�Q�W)����rR��:��Ѥ��Q>!�i,*�� ԙ�����?�w�Q`�,��rn��Lbj4tOcL�P>���?���渢y=�s�Y��6{�^����u�J��P��ixN�E%-����0 DT����|[X����WA�PnИ�˼o�Q.�^��퉰���t�����_��Y�K�}ĳ�#�e�5�,"o�_�AD�S�/�����%����	%��Ô��=���W}P��O�Ch��oFE1Ӻܓ-'e5��f������hG E����P���y�{e�N�R<��v7�c�?w6i�]���0���i�}���i>L"<w_�"�7��N�TN�Q�h�}��9��'�{�b��%��S'���D��ߗ\�1yX)�y������̊ǉx���?2���ꅏ3cE�4���d��%r��=��m	2n�2c%z��p�F���_�eLu��\r2wV�S���ƙ��}���,�	�Gkۻ�2�8��ϘR��n���P�������[��gs	�iK�uI΁�%�A��0&�F�]�YoD��G����!:���yIF�����p���ݍ�H��t�p�Sr�j�~)�q�l#Q�ơ[�A��S@GNXC�x��,�"#]H�\�T���[aRN�Z|v2A賂!�U3��r��Pj	{���9.�3���Mb�����@%���ħ�|�7u�yo=��.�@��T�4�HP�y$k����M�׵Л&�3�JW�Q��J'huy�W*�!^�ĩ�=Z�E(�J
��M3�"�͋I�Zmߨ��2W��72>@qJ�ޤ�e_&o���ndo���t�q�"��P´�y��������O'�߁~*&�w��K<:Π0��h"~��YT�UN<�OѪ.k#�Su�E���s�������Yצď��)���f��'t촄��|%6�\�(�Z6a��:��ԥP�˺��']� �G�2������'E�M!n���9�%�c�ԥ�/r�p�(2�C^�s�vokW��� �Xd��*CB�:]���Z��A�3�<bلͽ4	�+ۡ���i?���%����n�c��mҤ�����0����\�C�����X�r��D��|�="~���9P =��l���0�� J�?x�o+u����f���י�zɯJ<�l当��xe�{�$���HS:�i�-��)E�9l�3fI�D
v��W���{I��M��C��
p;㇎O�?O
��OEꖌ2�D1?v��$f��{�6��rD{S
D�����S�7+��u=�dU�i��'���׫����k�d���_�
[qK/-�Y�4=7�&��g�n�9�bw����jz�m�S��=�谓�h�{RM4d��Y��nSs��:D�G_Q����|��A �HW�*�؊�l"��V\���]��Kc�����9g��{J���e{�s��g�q[��[��_�r$~�~)B�����4(a:Io& ��g����u}��W�|Z�����J�6�Ӌ�6��xz�:q���N�%�a��4ח��Faw�~cK%]�D]6E�	��L�f�▷�]B��D�>��e�M��ҥ+�:Ҵ�[���s���=;�\П�Q�Q��B��@h2� �����I�OYk)#���/��ީᅩC��u�*v��;x��7͌!�c0��os"�D�jF��\U[�(�á�!ɋ��8���/�"���v���E@qaP�$�.ZW�3.�.�le�s�or�	��_W��|�%
"��Li�V����O{E7|�WG�Š�ʈ�P�P�*���="��-E켃=�e��s0hW�	�F�Q)ڷ���0�z!�,��~mf��-��n�8���~ ��`t�ً��fO/��\o�HoG�U5���qVǌ�,ܖ���0C�Ċ7�*Fh��}���/<��)�"���A_���,�0��:��G:�Cж��?�Tݰ:
��j<ث�{�ѱ��Z9���_�r= ��w�����IbТf}�ߠq˕�#:Ä.�а�Xk�Gq!;.�、DFA�i�������>V����(�Vy�D�Rl���T�Ƴ��,�#��a�q��BAڅ�
3�����U_B]�r���ͪ��9��p�����r��.,z���WA�ϩpQ��젔�]� �ZB?��u�"���a'��0f�*<�b��5�D{�9�Z)��!)� K��K�:�.q1o��n����;_c�H �[Y\��;���?YtI/��$���*,�w���6�:���G;����)V������"��[��L�.�ɀ��|�������f;���ݍ���X�.ロ	"s���/UxdTI\��"�i�8~��J�3
%�S5�NRC�p��7M��H��bQ[F;t֧E��s�%m͐ڕ���b�ޗ$v�9��;*E}��=������A���rz|{�����Y�N��ŕ�S��AC"��X�RL��^���Z�-�#�Ch:cK�����h�[��Z�A��,����h�D\��u�����8�4Z�7_v��T$r��Af}	�.���F..���WUX�����_��U�Ǆ? F���n�/���v�\􈕎f�C���)2Ð��b�ںn���R`�������4�.~��2H�kݑ}>����x;< ����΋��4:a�'DR�荐I��F�ɼ�rAcE�gO�o�hn�lZ�%�q!lʜ����ِ��M����W3��f�Z#MZ L�v�@����*:W[�/�h^�e�8����HU��ԕ��r�w�z��0���m�.�-� �L`�>sqQ|���.��y�Dq�sm�g7�o�,uŽ%-��"���~Q��+W��O�y,t=\S��=#��G}�!R)��h������;�	�D�
�o��_�����X����9���z�QE��O���������u��M�&�Kv\+�tn�����]�m��u2�`��ï�O��{-�6��
�BIT�,B���M�WyV����R�ը��N�����ֆ�l)�⻊�v�?�My�K���"�
U�
�MA�#aK����t{n�C�>^'$V� }����&��;�s;7;����ë�f���7?�u�zWa=�@ڨ69<�G�yv��8�8���-��� �H���ҙ����I�aU��DP�3uӝPo��ҴP��0|�&'a5�V#�Мk���y�U�}����!��J�)���Q�>� <t|��������������wlJ�^	`nCݓЃ�Qm)�74��S��7p�l���BK�R��l��%��DOn���^��#�Co-}����[���]�Z���A}��[��v$��n�����B�|� �3uV�qJNh��^ L�`oCg]I5��ż�L��w
O�l?g�C���Fo.B����0���J%?Pœ�4k��)0��x���ЄB��(J�;�\� PMɦ}&jez�6�M/��]â�DY r8��/M�j����L
��~q�3�A=�ׄ4�+�t
�f��'%.�J��@���.�?�/�?��t�(#��u�\��������.>��M�@��e�>T���2ᨳ�_/�֎<Η%�gNX�K��	?N�AY3e��8�Z $y�3��ʬx��9y�U���}��]xy�+P1}�r��J�i��	\K
UG���و�}i�7�Ź;�Z�}�B��1�A{LkdnngtH�i�l�/�B��>��m!��g]+��`ʡj\% ��s������h�~OkrD�@v8`J7�v2�T����sg������c|�����vaА@��.�q�(��pn�8�ⓨ�ش���e����]�=�����@��Q
W���
I0���I�H�ka	'_�BH�Ķ�pO@�m��L��W��cG�*}@)"Q���$+�T3�&)H�'��)^ �\HY�=�(g�b!H�e�l���>��X���t�c�07�L���3��w�m)�f�`3�8Rwf}Δ6�Z#��!�M�P�O����A,)�l���-)�$G�%X�����P��~��G-��$��I헞mT�9]�a"�A���w����n��D%���}P�A��Z`�Q�٣=��	�t/J�.Nv��M�'o�Z2�u{��l�g�+�Pc%�VA0�O#�XW�\q�3M2=�O8�js.D#soa����;^�X$�23 
��@Cz8�Íj�My���2F�]��)&�B�7>H�����4	�9K��m�Lq�����$O��`���+�ɸ��ѯ��
����!��x �[�̏�i�a��Z��іFyƧI�V��Z�ݒ����o��^>���W�cշ�f%�?]�������F�RTΥϵk��2uW���hp�))�����W��[h)��V<w.g�fCV^�VA�w{W��է�ơd��X���y����W��wM�D	��%D�ofqvj�Cdp����Mq�2)��޽cvȥ^����d�T�&��~�;_'���s���>�y2��i�	꿠"$5�!Ƥ�[�T٘e�ԫުY�Y�k����|�ȸ��/ k(l�t��æ�D[V�n��T�F��v�r:���L�%�������A�hPL{���a�jx�qZ|���Zch�<��v��916���!�A���]u�_����!v����B<��(��*G�Џ]�-��������(:#��'N�E�Y#7?C�@o�x�<ǖ��NdW���V��r:��W�����8���zY����?Ȅ��a�S$����9����)�����}�E�C���(�V����ˬ�;r��봢�j�{<��SDWǍO�F�����w�T�� ���5Ԣ�;�#:4��c�p�"������R��"v}�X���(�]���yB>��оey
~m��fAD/.Qz��^I{ Zіsē[�,}��?ָŃ)�����1Wk�����@�}��n�/�PA%����*�Ŗ�^�e�Вo�����nCe2���J'�G�P{���ϰ����5�.��w�ڏ��x|��cS�����?{P����/ZS������s�u{*�b�j�� c���t�/�ʹ���,i�|���V�g�R�2$�/��T���gs�n+�L#�ۍ�-|�zV&k̓�E��� ��N�����=����9��9ϐFǨDzQtM��}YzO.+��v�����'b�W���b$��I��zɻ	7o�X����?��c��1�c�+}uy��:�a(���r���f6�yj��k�B�t@:*���T��q���@0����؝Z�#v��r��Y¯@�|}�v���n��}.k�p$��4�B�F�Y'�-�A4'��0���^���]ڢ.Y^H`��uW��`"���	��4�๐w��G7|_����6[f��A���-7������ίT5�ލ���b8VKJ��O�N����qE�+;�F���H���͆Y��]kљ�H�q��ك@��a��:sκ/N�)f��Hzn�uV��Eu[�Qc6jz��$�Dy���Lx�$�YUvo��ʎu�v5��vEp� P�<E�עOh�3��EI!����c�U˗��i�����
�>d��}vQ�)?��=|�q+r�ْ�������ȏ���zgm�N���w$� IT�Ȟ�gX��AU%2�
u3l�b�:�;5��xB5���\DÎ�\��8R��X{�ɀ����_�q�I��F��w[>p:e���k��Ѻ��,2Gސ�����!&0�,�ɮ��@{�$��E1"YG�/����*S�W��*�5)Oߝ�*�,����k$;L/2����j$~��M#~+�MC4�� P$��Oz�'I�q
�ǉm����!k��[�����^a�cD�:ڢh�89a�l<���$�\x�NF�~����!������j�Hl��̡�5h�cci.���]&��v����]��QG��[o�(�FL=I$J̊A�6N�[&a˗=��F1r�?2�,nB,��	��8�Z�k�𕁟�����������֍�R��Œ���A�|Y�fAhh�K����G���!�@�1ي��D��$�p����@p�!_FaC�i
��g�᪪ڳ��#eX�*�Vcr;�0N%)h�n���(����O`E���vu���s�[+p���hV΍�;�,$&T�[���mlFp�M��9���E5�?1��C6FVň���8��r߿G�=>�D�d;�șc��SKM� n~ �}ﲖ-�1�W*PQ㦂�b�d�fB��`�T�M���E[���_-jO��lc��rW�Q�h�n�T�%��?�A��H��#��E�7��"�Ks���cbj�ǀW	�{��t&�{�t���p'��}�'��#<���tW�/�OGdo2�Z�x#�S�-"�v�H�@�cM��rok�#ꋦY!��X*�`����ó�t��6'Uh�n�%.�Z����2�M���Я�38���Y�г"�;&���.��s'��2l�b�Zo�ć�@w��좉�*�\�g�z㹄�����y����`��Ȓ�~������?S���s��15��EDw\�Xm���zl�G�"uf~b�}�3�G�6�x�>ћ1(-��6%�D�#㠐?֕[�
�/n����������i��9}6�˫8���������	}�ӷ=9Qo}��{%ٳ�^�>1��m����˳,�:;y\���-BV9a$~�R]J������\N W.�BO�l����:k��=t�Fii���O��s<n���.�љ��~[�8��W1�K�.�)U'���p�b�,�m�|AD�*V3�ńfqQ�N��ǰ��q�q��T�ƙ0�n�L?oh����ӣub	��RS´�[�����TCnx���c%���0D.�
�{�Ғ��˥C�[�����U��M��!�"ځ��~�g����h[��`U�YnIk���� ���ydj+��]c�I����QR�[��1��e���`i����X'?��}���O�e��ʘ]u��B�sk D�-���ˁyx�̟�z  �u��?Ds<C�+�� FP�Ҧ�j/�wh�3���w�LD��z�-v�h��y�r$�=#��9t��g��݌�e{�_�71ޫ�x4;o��]�0���Xg�"Y	g�9��mr!� :��/^�ǃC��{�м�{o�'�x~ b��<7�ǒ��n��Q���2J�䮰�XHg��K�b�������0u^�[n)�l�uF����zMg%.Is��c*����*���oDޟD�.o{R��̀��s,۬�#��L�P����]���r� _UL֭`0v�;_�d, _��Zv�_�%}��h^���*ꄊ��
V��2-�ؽ_� �,F/55��IkԌ�"/�g�<Xi<c�e~w�_�?Ym}��Kq�^�E#X�=������-�2���g	?���+�t��d�ў�9��#��7٠����_X5��G(��3�d�]$|X�ۍ&�E=�e9�ЛFgT����ϫ(S`���qFY�J9�� ���w��;%"��� (��/�)H��@]�lɍ�tp]� �0�M9-).�y:z�&$��*�"�cS����V�$��2�yu�!����2/w#:Ւд��rr
p��i�>JN�Pb�x��c��Nү�����5��{��M��)!g{zc�#f�Aj	�_.��H�M��+���"�}�W;�١M��I��j{��V["�k�lQŌ��&X�� j� ���,>)�6��"��zw�`{���9���:'����:*��ڹ���[�V�i��Tׅ�X��=��d���:��(\�5��L?�D��U͔�h�������ir)�E���	'H��>Iv�m'��@�$ʚ6�p���9&�h�ms+'S�"���Bo<��l�kuW�g�^gLw�ƀM���3DL�[4��xY?m�9����uP~r	�2��u���XN>�����'$��^��@�T�n{��b�N�]ܨ��I�*�h_�_� .9�g"����?@l�,l�f^�%lx���$"|�k�0���5��`P���}?���4S:�؏�_�\�[fL�/������2]�)Gy�� �f�����c��a]��p�d��0IfC���aml�1ε�w"ʶ��6�4�bC��[��F^q�7������$�_P%��a��\e�d�9�a���S�-���B��^I��z�`>���ό��U�����nMٜ0�R+�$񕹟Y$��"�E ��V�y���#����6I�>)�v=�YkF�R�4l�׹Ԝ?`��k����?�nG8�FN��!��[4`��[æ��9������-5�%�rD���:p�KaG2����XߡK�D�K%(a��pE�,�	�k�����:!-��ep��oc8�%�ѧGOڍ^"
�`QCf��3(j2��~�������+�'�s��y&CO[L�;jQ�EC�_n=�H�w�wt(R�'C��!O�BT���)�ܲ2�6O@�3�o�����_e�L)*�P�0����#��/M��`��7�ʮAQ���z�!�����;d��k�x���U��{Т��$m_j#�	>�C��۱�@�]���]��a��q���fx
ɷI���A��`o�0�e�3*Wz?Gg���֋[�b�z:rřǨv��̬�(�5D�%%˹G�� l~�\��^u8�{"�M���s%����k9��'v&�7�"��V�+/�ϲ���KO	���HV^�QŠHpc�X����		GG�%*N����9�Fd��(m?ms�U��nF��n3�Z�&�� ��<Σ#	�}	���xga���#��&��"�Aj��{jmضj��4��0y1.ßqn���n�����>7���(vƨ�p�O�w,�#,-����/��*O��te���ȶ�}�>q>Mur�ͣ�'�⚶Q�e<;��a�%����������h�5E��q�h�JLb�1�<!1f >�cﴷWxf�����b5yZE�P��H�N*D�����[�D-�?��1���m���/��gtB��%�b~z�"Ηr�O�w��
�鎾M�W�
�;4�&C^̛��'_f*=Vl��b'xSi���yU �/L>��r�����0C�k�˦ےb!_��ƌj��k��zJ�cY���;�B���9�����7�s�(�Ⱥ��4y(-ޙ��M �U.��Ԑ�����9��+^��V�(�q�^�/����e�e�_�'��^_tiCρ�=�'o�f AO�&#q�0zL��-{{a�������V�kQ���F�ZnG���?eN]�g����7����#��&Kn���`�����qt����.�
��1�՜1�.���+����Jญ���|�g$������~$�?����k�>���jַ����:��Ӻ�Ik7~Y�_�n�nl�����m�Q"��;�A�7�'�z���Ap���g��|S1�\�:_�x،F�?֕�:�XMYӮC��03�A<�6j	���\�ܷu&@O���;�����E��H��23�s(��/ԭU%$�R[�T�!�W w������Q�=������h�*BԸ�B,��.���� +��.�L�]2�j���:�j����CeCV2Oa!~o��q/^���9a��_I>����Z+�! ������f����JZ8ր��;����BZз��r�e�����[5c���(�2�j�m|�.����:$�sMt�":�s )]1�*��PCܑ;W��G�G���a�dU0�W,(�������Ѡ�-�u�g#��(�Èn�ɓƈ��D3�ܞ]�J��igD�IZ@�3�+�|�c�]�h�~:F�s����/�P���:�k~ � ���{�5:_"��N+� vq��.�W3�� ��@�6�Ex.$M��.J�gݞ��,����)Z䥉 2�ɼwz�s��Q{�̨�{����w����4��ӷ\���ƅ����򅓚T�`��U�=�|k�.^�c�k��<�K@QXk�-|�����g��.M7`����I�x�DU��R><r{{��o�{8<�>a�c	(�q2������v���%�2�it�N�T������
W��ޑ�5��?�� ǐOه!�J��z���Y= �*�zОT��������s��e>�O���L��q��x�o<�Z�.M_9�r��^rr(#�˻g�3{z���5��-6wch�B*Fd�	��v�Z4C���ضӑt*��X��˄��Ed��ؓI�7�ee��l�!Aq�/�J�aD�iʕ6;���Y2�f_hU�Hz�9@�q����7�΢H��]��ӏj:Ɲ������w��Y��c[�;�?C��^������L�$?mi�Z�;TwX�\�<�K�2� ���?�T���=�f���ιv>�A�n�ī��s�/E�8�nRDa|��i�����ΧLDZΦ���杫�>��_2�7��������5\�fFP�iD&�xO�d��^��VW#�Z]\5�1�z}7�Kä�:�Ї¼h��*Ē9��!n��+܇UX�7g&�?f"2ӑ��qz���a��S�02e$�sR�ف�
�r�r��Mw��������Ǌ������Eڅ���]m}�����!ӎ�g��!����P�b@5���UN��,�Z�N�r��(@���}���J�VloC<� ņ�J��j-�aavJ�.���������5F�X�� �l+�]��R_��u�,1�PǛJH�X�T�.�v�W�;k5�u9�ka�nZG�����o�86�ɬmۙ#%.��!��zU6���������|ҡLm��pk�4o3١�	Q��_5���1,�amXˇD���{�������E�-h����j�sش5�k����CR�c@/&�cZ��d#���f�&��ǎ�e1s���t�������)��j�z�MS&#(��V.	u�5G��Cc�s_���.D@��,(�,#U����(T�I��8�b�W���IBb���d�.e/?�>Q��S�$�ot���.&�r��(.�R�����<K(�G�"���㲛�n��έ
�*��[��n�b�E����������[1�T�+��7Sύ�S��8@w���Q�ҝ�#^C����?w$��ԕS�5�9p(�\X��>����rU�|��gh�8�[��-$�"��U�;�n�޴���d�L���`��D�b��$���g}�d��h}Oȓ:��qp5��l�����"��)�3����9����*鎿��ގ�Mdnj�H }H�f)�m�w��xd�ޢ�bw�i�Y�_3VA9h��ϵ�sӸ`��*j=%�U V��I�1c��|E��#�n0����{X�d)�NYs�=,K��k�s>C�l��v�ngkQi����c	�ۮ-z�U�3�r9��ܕ��{с>}�����cyJ�~F�<�.^��P�sڏ�49V�b� @��[I��/�}�*��N�s���H�7Ɇ`�*{l��[>eW��r��o�4*c�^u��:6*be�u��d���I��H'Wm5���Q�$�PZ4�Y�ט� \@V4��nߧ�G�1�� -�F���z9]��������@����O$�1����'t*��F����ʨ%CAU|����D�ns��0��l.�U|������������{ּu���#�YS�*����2���%%�O��Q���Ò���J�#�c��$ߺ��etXf���p�-�@T_�N���;��ٍ�����+&TC�k��~|���Y�[� I�P�Ai4�a_�<#�q2�f@(�����#�S��Ȅ�r/*���/r%2�>xٌ�r���>��|r1T�>�B��|)��)�B��;�����k': \&ŉ	�́�<pb���Zc��}���A�Dԙ�ݶ	��}�a�]���AF�r���NJL}��o�5��3�l��Q*-ݝs��;��T�
�}jd����H��,���orx��t�zS}_��u�u�KIԯu�>	���(�6���r���ve$y3$���oʫ�騇�� ��=�N��9۽h���"zWЭg,-B���r*��� R"���l��ig9Х�B�]L'�܋��nh1��_�"�xo:O���)2bʝ��ujB�m-C`��� �{k�9�3�G7Y�p]�^�;�C��c�M��V�3d�'.�H�|0H%��n[�6��WR���	gh�cVBD|����o7��;W��~�&G��_=u��4@����^g�1:��`�?§�n�o����j��}R�r͇����3����p��N�|7�������7Jݠ�q���Ih}Tu�o�����|=���}{`ϼ�iU�k#�I%�rWy;��6IZ�����,N���⢮gv/��A�~���O@�E(�i'8띏Ɂ�˯c�T��I��.L�2o���(7�ǚn�臌	�2��2�Xbv+���Rg����!tI`�n��/�/s�xh�튻|�J�a�kBԣ��*_�� @
^��i����4w߽�<�b�V'Qf�5����-���bD����ɲ([�)�����,�f�B.
����=����rݵ0��46G+�X����Y8��[����:�
'�iH����	���E����ɨ���n��V7+��{��"e]�i�n`�:F���ǫKw�'�B+�U\6^Z'F>·���P�|t��p=�����Ï�@):]��g�)�U��ir�߷h�iB��\�"=��D���"�L>���RZzT����k����Qn)"o�a���&}�) Z�
6���:gʩ+�_@>�S> 6��FMĲm�L:|J҅���G^�}�M\^\+/�"s[�.����!����,�4�j�i?����娣1�_�r��e伤�8� �$�UT�<\��B�wcA��qd��2=l�jJD���3��C��]xQF�����*�[^��6��Y�}^�|�u���[b���s2�g�(�!����V��(�D�{G��8�ȸ���/�7j�Y�c��*�Z��o쎃V�I/9�dp�H��@�Џ�~^��#�=b7��^�-�<�\ ���S-WMX@��
}3Ŝ",�TW�A	��k���x�́�1�4UηX���ۅ���/�W��b4��+H�
�a�웺:\���k�܂>�o=�)8��Ci��
A@@G����2� b��c�z|*�"Ъ�������1-k���-#�Q�m���d��J�����5��)̶���O��߆��_�G�:t5x,-�'y�؍=�'�v���&�8���(��p�ҳ�@�qGQ�F!��������Y7�C��O!]��x�b5��+�&$��������O��+�(�Ȩh
EJ��D=1�����R�N�i�X��/k��̫�U8 ��,�������-EM������v0��1bF��S��7�58.�av,faŘ��^��"���u�V2F]
�H�~-�BH
���0ַU�Njps����I瑣���j ��z�^�N��v'����F/N2B�<}\�y$����z���Jm|g;�9՜I���Y�N�XE� �2rb��(ȭ��2U��4�Q��3J��cԺ�|����?g»J�(�����mVZ7���h���s!UlD�,�~+-��	8���a�����/ٙK���&(ǳ���$v��0������!Oζ��ծ��l+�<]�+g�R�?��J�'���,]�3�K{ţ�9�e��+#x��t�?f]�j�.�26�� �E��:C���=�~C����oN�H~-V5�$g�a������r�֊:}nf"������!���ٙ� 	0���� ���Y�]݆���b]7����u�ֽ1�i?��U��@����m�o�������N4�qa݈"�U�>H�����1�xc����^!�����a+s���/o|����3�����-�����+i��:Ǥ�U�S<��W%�0�����O��q�3��(dQ��2~�;%�Da/�^B��� =�Ed�s�V���a��R!�psE��$څ\�s�%��:Y>3�J � -����eG��;�'�d4�ʼVۺI�P%ė��)����Ƿ�c܄��7�c�F��wK*4�Y_���1M$���Aj$��/�9�J�4��!���N��) �)����u<�N�$)wW�K� ��1B��6�>mb94�9Q�·���2��>t�%�~�C�M2�y�`�~�)͞@$�}4�Ί?"��Z�:����6�:r�GV�֛��2��k�?��	K�&���EڱX1�5��Z1�[�~e�\~���kv��m�4�a7-K6{zgl�ū�G���S�:����`�)
)V��B��&��3�0���G#3�5�N�]��`ST�E�}IҴ�(�Y$��Fቈ�~���3hTC����a^��O�Qcѱ �ch,����4�'m%�E��|���>H�(',��a��� ��y�9��B"�d�X7"'� ���z��D���n.oq{U�xw>q�Q^nٙZ��C��B�Cj
6���x}@�|��:f�z�3�0¢���r�9�3�V���{�#tM�棸^N��x�s�ZS���4������w�!�DE���[�sjAI�����i�iOY�gPpF]�U��$0�+�T�8�W���y�'k�/�!�'�n��J���: EՄ�����<���/uW��F(2 lw΂���5RE��.Q�&C�
p� ����h��2���9���E5�l�{�ynn51�ޟ�0On�m�OS��Ā��6�Y�Hq�=�ǣG���ma"8j�pIzUX6	,�V�o�3���0���r(���Z_!���a<%���I���a����eo*#�?dꈟ����0*H���	[/4�ʓ�T����o،A@V�3�6}��4�ݠ��qFaO���6�}3:���|Jm�n�3(�6����^ ��Ť�jKU���F�os,����6��"L��'�Ls��>}�I�?�394�����6�d�NE,k���1Y���}C,���Kk|���Z+>|z�H	2T'�Q���79��ȷ�֔�&}��d�� ܾ�'͍�bs���RUYu����G��K!2�\�i��Ʒ��ǃY��䐓[ �k����?҈���{w���`W��O (�d���J�|����L�<2�P����b��`t_'���G�	~��O%Y_)������s@�FMA�0C/���Ús�\J|���*�l+V|�o�k^�R:|~�I��4N�9�K`�,�C;tm���,�^)(�e�tA�(��c3��t�j1/Hk�A�q�)Go&vW�d���xx�nm��=6r����G���qr��K���,��GjE��?h�y��/hX"7�L+��VP�G�L�e͖� xcd�b�t���Мb�>�x��2.�G�_*{��*��	c���
�t�.���$*	W���h��uHƚ^ӿ�
.�YNb�H�N��Zl�d8�J҃�5)�8����Lb7_��m"����SxI��l��"�o���ɤ�4� ���7M;�]7�����	t�1�A.Ea�6�ߘ�����{N��~2[���{�����#�wEI:�r*R���(��Ik�:-� �i����~��"j���`0���f�Ak�H��Ь��v�.�a{�uS���_$��ݻ����o�I�_ܗ(>,�w�)"!&	��C[H;�Ev*��L�f�:$�~��&�`/e�{q�nxT�hV�<m�CVu��"�B�4=Y���Vi?��bw��%P~���ep�ߢ��Ԏrj3�d��BiBf:�;W5Bk}�g��#i��A�v�������ʽ��?j�{�@�)h��]�X�����CPY��g�5�ɳ%�5�1���v��}�EY�C>�`��:6e1�-6�D4�lI��W�@�'Ԝ�ҕ�H6��d�o�}T7¾/c%l@��ӐA���B�b�L<L˪�v2VQ;+�ʯ�[��=��xx�c~���q������]��
�[�%��*�M�)p�:��mE�EnNW�~"m����˅�I�@(^��9}��@W�ɚw�3IH4�3�O,^{���ý�w�<e�%}.�.��6��y���;��P�	fz�J�OY_j�`�sŉᾎ�ƕ���>IL�t1�l��1˫iD�e[��pZ@2[ @������ں����]i��k>o���Ȼ�����&W�
J��`^�x
b#�+���#�ב
�6� :
錎K>��d(��Y~Ň�1�P2yz>33����0�;>yr�����x1?�� �f	Qv�����2vJ���ek}fb8g�i����1_��E�Kl��`ғ{�gF��$���S��y>�H�	����%)=�>cx?qX����p��� ������<Ig>c���D��V�	ߤ;j�PB�a��\������^�qb16wc��Ҧ<½J ��9�ڳ���u����@.W��VR�Q�-���F;�H���Ax����V��0�O����8BH�����㴱!G���{��!*	�{����ѭ&���H���k�U��b�m��/;@Vm�g�\@Ķt}
��9�L���U[~��e?�_�����2"�x��BW�u�������C �~Y�O%�>+X��k=��
�$϶�up�˼�m��tB%p��P@�9���$�nF��/�`�:��;]��;̇%���;Ъ׵Zh�������*�+5��j��jDc�P��NU���Y@���lB]OS��$�\��s�L×X�(��|e���;�Q����C�T�B��?G����(�ē�7�����7�����+��b��g�
@�b��J��N:(�)i=��I0���jő����ݯ����ҹ������^��{	w>���������-T5���§��Ê�rm�##ĺdpP�*�I��-q�rE��S�[g�5���3�"?�'��թP��@ꓫk#�j;��Μ�_T54M�% ����=a1�����t;'*z�\��[�og��F�֊~K<ôJ��$�@)��#v/�{�5�	�U�E��yMЅ9�*�MFUwߠRz�������qr]Y���т�q ��`�i�o��q�0_��SO�Ýc�\�|+_PƙKM�<��3k�q�(=�N����U�����b=gI�)�?Ť���G�,�;@�á�z���@k�8x��A��/*N+�S~l[-;x��"#L��u/F����;�䝯�h=p�w�F>�q$����	Ғ����N`q�B��Й���A����	R J,+]�3�ָ��{v|F�[���k�~cu�r��>���9+ ����[@�!E�D�5�8�ї��9���[d&9����׉;7=�|��B*Hw8�A��E�8�+�ο'P��ٯ��Vg3W4���<n��Rg^�,b�5�¿���@��A�;�0UH�{%��H)�_,�vjJX�?|�b'*1��믓�s:����}�M�=�>�� ��[s�.��t0�ļ��� �ɛ8X1���0�5�7(�?2 y��AD�����R�N�	j �έ4x�ǊK�m���a��"V�ZHQ�v?b�����QKssm���ݞD邏P�~RH���V�:�sf{(H�����ZsI攣�J�c~��>:m�#S�=�e�H��sb����Ɖjd����+�$�"���g�����و�2�\��l������W�>U=��u�{���L퉆�q���
-2i�I��]ıԪ^~����i��;���m������Zw܌&B��YT�A�y؂�U2�4��@X �(:�րi�"9A��K��\j:K���C0�7r�96�z3+���H;�Z1�9kRLm!�Qp�^����p۷H9��T�w�Ϸ�z�5(m+��yv0>���'���ҿx�:��Y`s�����H�[�l��
��;�q��E"��jGk���0A�Ǟ���:ԓ,9�OUb���ɘRB�L����<!M:0�k��N)��1$�6iF�IW���"�ӷ6���h\�j�J	a���Eo��w�X��A�`��>�G�)�j���x͜�����#=�b �� $uw�Z�X�]`]5�]���ÿ��s�,5�Yj��B����Z��ŇxQ�O�<�5�w�)+�Ze6��%D?�i�i.�`�5̄Yy"� 8��,n(`0�����|�9����f�Cb��㐅7s�n�݃y4�YL��zH^��ث�}Ew]O>����������\��$G}��yԒ�g{`-0*���`��U��Q����B���מٲ.\�W�T#H���.`�;O|�Q=L����<�������֨���!^�R�����T�Nb� fI�\�)mI��ĭ�NF�֗A�z���k�?v�o�Eՠ�A���-�9y]���;BM���E��ZJw7��v�����ƿ��/��~�yH��/z�v1h1���Xf�;O�4]��Q~U��ܿ=��.Qm�x2s��q���R*�cv�szy�S!��gv�;� '�Q�Al7�#2qO��ӽ!G�@�G�ꍤF���^�gG�[�7ky>����'N�{_`��*����;P���^*��mɾ�%XH�e<�WWE0F����W9���7ל�mj�@�w��1�:F��B	Y����0���ѡ����M�X.�е����w�[�����4��/ai�����4���G� �Ȼd���:@ bA�<܆��@���K��b�s#���1v~n��xVp����6A��x)�Xmbw��fo#�%��w5���J��1蔬n~5�Up��:���i��֪�(Ir;aBgU�R��`��%�6��[G{g��5'ue�.�-�l!�l,0`������$k�w�+u����\٫&��\U�&dA���h:���C4��u�)�S�j3�E,�8r�,Xb�uh&^�:J�r3|��Ɋ(��6Å�����Z�VQy�Qk�C��u��G�����F@miŐ4������?+�� �R0�������iӐ��K�e��E����B�a�+�Z؁�׎����~6��8nR]��N��n�)C4�Vtv~�cY�J1,�Q7�sՂ�y�1����+���i��+
�q��:V����2�bw�R�!F]x��Q�rJ�>��*��}�:<�8 ��Q?\�~���)t
��l%�B����u�T�v�=Z3�3���Ӏ!�U�
�JNm��R\يE��ۏY��m\�e��9�f:=sV�
�j��@��$��N�}�چ�����Q�(���n�<[W�j-pg~G59��c���������ecǵx���/�oG��R,��i�ce�H3~����i"G��uW\�:AM�H�>��X<�_��+�n����8�;����E���X��j��vInƛ*�hc������Z�~`���bs���z6r��E��B�ʅk/e$W��{��;k���(���㳓'v��Wj�׸���0�N(Ѫ�aΨd�7ܔJ+��"//f���%w�%�����H��3�b�]�"��Y:F�.{�sI1r��Tq{�ٙB�Q���hĊ�J��q:�F�#�}}c[Ub`x�X�\��cةfE�"F��M�`]8.�w�ũ���s1	|{ٖw%~�$8RA��t�� �	ӱ�D9��h�md��H�H9�fZ��������A��d<�9�V/ЯZ*^(����'���6aTi,�,d�r�Cg�7����Įt�%�D�`2��Kx� �t��Ψ<O���/z�k7�T0�6����	�N��kPٵ[�-N����ވ(yvb\�e��`ƻlץY���:�XA��e-`H��٫�@BM��W_Sv ���<�n;�z��DU?i-�TZf��p�y�R��G�)�d��[x��';!�=x��h���fn���Z�PC�K�љ6�OP�WO]�-)3/��R"�XF�y�U.�ar%�L�˛H��{��i1�>�j�9�=����]�Ag��x���P��~�fhb̰�<�0��{�;�!	Pd��*�EX���*4�Vߦ �+�:U��mw�%��jf~6oi����^#�t#�V���Yk���5b��!�^[�;�F��i�a�"Fzz�1<ܴD!Rkk��j=���1U�[ ,�	8��ͬ#�x� b���d֜�]�S�=AFAF���O�u
��"]�O*3fV�:��}���zx6�O�p��s��qD��P-��D��]�歉��
� ����N�~���>̒{/�j��3U�����ew�:%F]5��˜��S�A�����N&tt9��80�do��o�MKE;f�?�3�'KdT:
����=��O[��
�KQ	�����=��$^�������
�߼d� C$܂2�	W�U��=G��\t�5~�3�?�L��v�j��x�u<�sN���?�+� �ɻ�k@�!��&y����:�Y�[��xH����
���O7��~j���H�Y�D֍��,���N���29�u� [lKm_M��*,�nU�睻ځ�qL��.����Z/Y��p�-h�R��w�_����[*�&p�MO����"����iN�������J)�:{�~�U�bTl�g�F1D���,�H�������0nu&WE�iYi��>'�y�s�j6�������J�Y�m'��d�y�x��5j��12\ M	��:��9�^��qH�'�3'�8;0����륅�޲lɑ�p�}8��{�~]�H G�~'�ɑ�H׊��h�K&��hЌ�	��i�;���[�3�dr��TQ-�am*�k�P��0�$�vo�I>:��_���֏S�(�Cﾦ=�ң�Y�r�����v%��rꅧ�f�ߙ�� �}]a5Rp��]D�����H� :j���Z����8���Lb�\�>����	Sv���%}<֍��́��Rk}���m�Wޡks!�0ſ�_T�h��vTSN�6�Ƴ��S���T���B�
�UB���u�l��}��#q�z/a�ac���u~HwY'���>F�<�szk�����I/s?�Ö�,����gu<�()�d��
n�x�|?����,!.�pe'�9ACOh�kZ\w0{v�wT<�Zw
RX��Q�|	��ג������H{b�>�~Bi/n6GX�(!It�lwo�G�|a�ϦH-����{�>�F��%n(�{�"!o<s#`�$[xqif@��Z�x��3X��u���Q���k/�^9���y:I�Sg��@��zLBDhЍ�w�[d��"ı`�SE�T(�����'���{ఢ�5��*���X�5� �Mݶz��w/;`J�T���#�S6_����6�_�S������z�Q^��f��G��ƜT6�ס4��W�~����p��[��	�ǟ�|�m0�$Ix�Q�b_���G:�����Wra����􁳦B�jUv?���7� ���su.T�d�iy�A�0�V�}v���@�}P�� �F�(�?�!v���BE�d���2�+V��]\���ٹ��T�{�j�n��H,�����_X/|>�?0n �X囮����o�v@Q�aH���	gF�FHo�-IcR�M����z��@�H�kt�c0����nJ=�H���M�9��� �5(p{hX����!����A�Z#��H#Y���͔�|Ϫ9����qv��Ymx���p�ӡ�x�'x$w$y��_�ߊ�ϳ*Ur 6��4�˝�r>���J�x�� �$�v����������tj\�BD�aj�.uX��G�iB���m�@exB����j�ۄ����m�sC��ca0�'-q�o� [f66��j��ib���:"�/��:��$�$�mW�E���lO��ڊ��S����Y�c����M��?xz
�)���|xk�h��8��\���$[�rr�{bD������p�#��b
*�������.<}ܥ'Z�Y����v-�J\��Nl�F���[*�@C���b�g��B�l�1���f���gk1�\ʲ]��Y��zȓ�1�������	�]Lf�Q
��l��9�n�K��:|QoğC864?�u���HzT�p�g&�z��ɦ{�g�>˰%�	���Lk۞�k�5��q��[^)�.w�����t^[�s��g��F�����2-{��"!��%j2���K��r'�����o��rq0���+�6��}ސk�[��up1��S����@6WB>Z�v]��t�m-E�d�ШR��H*u؊�.6y&���E�����]��m`���G�]l�H�O���h��*��;F�0c���Uj�p�H�� ݃�A���fZg���S���q ���va�2)�?�M�P���٥X	I���]�"���m�{�,�����X��@�j�G�v�Ǟ�$k 5�7f��Y����i�b�7t�����l
%(܍2�V�>��,K�Q�J8�J�+/7%;&05��b���#�h��Щ�|P����t�f~���������y-8��s�N��Dk$`�b�z�8G�G��(�Z��B����*MI��.yW{'�`7�:!D�]�OM?o�A&��!�&	�����HJ�A��.g��?��3�C��l%l�F�;F���j���c�����{���b֚p����ʈW2�ds�һI��D69�D�GN+���v�u��u8��SP�1�#��)�Ț<k�.�4�MuMu&����
+�1K����KCc<g��4>�lV^o�s�>t�p���BX�L=ۦ�:_V���|�&x�o�\��У~�r7�؜��[$��/Y~�,O�)68��%j�PO�d��2�5�V���C%��p�=������.��s!�P��w`#��yCidŁ��k�D2$I�FM�j��la����0���<�e�j14�-[�fJ���[`�K�-�۞��o&�T��v?��}��},�5��k�꽂�YԸ"�������q����y:�x<Ǳ��A�
���o�b�C�ز}�����8�G��7��� Pil�cDZ~���3����= �F�M�OeV��3�#�����7�#(ƅ��b? s�[+f�����l�P:��&�3�֖��M�F��x�a���nǊx>�V�&����m��N�͹��L�X|[� �F�Y��s�i�/Xtt��_i�Py�A����}�73j0S:������#��=����h�� 3��R�����B��ٻ1�9�C�i���?�TQ �EЪ�A��Bվ+��$ǀ�j�*N+9A��Oz*�u�t�ɥ��]Y����I��+�;COn��t�pp`�@��6����f`z��I8�K5��zꉍ�_�k���f5zc��h�
zt��S|r/z��e@WL�;��s}�L~�ۉDP�1�6�9��]�!�g�O�ۖg�����2�L�AOm+�e"��|�й5s۫��W!���q��DQxL��+r鿦0bp���pe�-�[av�t)�Q�^�w3
V�����Q�Т%M�&�W��-�*mf��Wh�"2-E����}Ae�&����G�hr�5�	���6��,`PD+���ϥ���,-2�Y�B�[�D#\@;�C�Z-��u�^�=+�=��j�Om���!��q��S%�2����;� Ǣ}4nY�(\<���Ł2�g��]�G�M�?]ֳ��P�<�
���n`Cv��E$ݰ����vw[���
����G���{M��M�%��&�\�Oz��l94f����,_��`����}�+�6�D��[e�r�0�|W�w�F��"#P���_�nV�vs��.������w��c߿}G=�%��pt(����D��Q��k�(�>��ψ<ْ7Io)?��n���Y�~�bL���D#H�#l3��Ra�t��p�[�'P,�5�Et� �r~B��Qu��'����K�8�R�js�M��a7����f�:�855[�L9Yd^���3��K�_g+$�wM�"��.�.D��5���)���2W�T��I�3(h+/�%a�=��w���~��sHϒI?p��{y1>%m��M	�o�`�sϸv�Lp֋�p\o���Y6�9,���e��hz��!�G�.���<BOn��O��t���������O����m/�@������D.XA�8a���2��ni	TG�ݒ�ns&��c_Y�_%�G��5G�#�n����)��f�0-θ.�X�߯��C�+��f��r�;�-����0�M�w(�
&q�VA�6)��p��B87N�|���%~J����hEq��O��0�8|Z\6U���[��>A<��\B)�����jHR��S)�󀭋�@2�-�ww�|
V%I�;*F0R���f�ء^;��Ӕ�[Q�h�#�@[������:i�M��vW��8�1���T�<��k!��l�z]�m��=_b�K��߯��`�	�:��}�M\x�(%�%F�ụzѹ#�|�Yɢ��ey��\;ė�(S��2?R���'h1�1%`��?;�^[��JkZve̽'@���8�NQ&���Y�cQo���l��"[������E&O ���bj�-N>y���y�P��`EM"�cc�2zj���-���X3�^��^�^'5+�� �*�B
;+G�N�r����ۓ���;Q���(�4E�v�^ ���T��m��2������R�u&M5 �B�Ȳ��O/��=��ߤ(��ٷuf� ٲ��`<��</S�lm��k�fq����#.KI�%�r~���R�s���h�����7�7��}*��m���l֭�1z
� �9��甑?��A�IªR�7���;�MG�	$�py���Im��L����1�Đq��Ռy1����@H�mE�+\[S�p�t�ya��D�FtN��(5�U0���(����G����$]C�)���MN,&�ъv�o� �E��T6�:ȁ�k0?�(� ��G��ԖM����y�9`{����s,L�a���W����Z*tX!�2(��"fuc�ds韖�劎�ǁ]GX<�Ll%�~�B��"�x6$CkzO}�0r�>��<!�V_����L�%��'��ᓏ������[A�}ba�	��$y+�b�k�eLy15\�|8/�xx@��[G���\�{��l�*w���%�v�`�vN|
#����~d�|�{���vz�.|:G��yBPu=I�4��`��pM��ؿ`�}���|39�kV	`���{�0�4�G�y�k��˒��J�gC��/ܿ�b��f嚁������
����9��Յ�D�\h�E}X�k�����o9}�h���v���1�0�Cz�J\@ZA�l]q��z7b����%�!}e�B��[�G���Ü[��BTy*6R����/�e��9�#Udk�{�v�
6�45t��c��?s ,8IiB�S�7NWk�(_k��$�$�]y�z r��G �>�X��[�1�	h��+B1^pC�t��|�A��(j��|�k<�)6-��V��"��QG�[7�Vb��@ �l�]�#�]
��<d*��`&������I�f�S�}C ��4�����Ueq%������>�n���xZ�����|o�O})8%Kk��q�he�t��szZ5�L��!�?�$z�nc΍�LM�W���7�hS�E��-%��ڞ4�qӇ�~"��o���stz:؛$�׏�>��kp5��0Ka� �Dj�ɗR�Ou����������Z�8��jE8�[�/�~��h��4R�	缚��Ϛ6��74"��<{J� ��gL$�C�Bȥ Ҿ�W ���}���g�H}�hx�} �y'�rE�6����
	)�^=Ƃ�٣G�ud���[�����ɿ'���%-�n�ɍ���xy�d� �М�� �5�_m��&�Z8i ����G��5ډ�|�0�\��)�3K���P}��?�]z3�����:3X��M��̿|�{H
���O���X�r+�{d��C���߽j�#xPZ8s���	o����1+C9�k[���~���U �ł��G���A���Y�yj/�h�3�\�&��˨"u�w��ph�q���!���O�z��ն,V�����J8�:�F�_�V(�T�nmoL;/䨢xU�#c_K���.�r�=���m�T��\�����U�=�1jo���B.d��Ζ!t`6��#��3(��8t]��[�qu����\�L�YB�}=i�:��y�r�0L�߰Vs�ب�?��{h�lO�>,U*N��eM�}�d���FV)�P值D�B�[z{��n��z&z�$ާ���ٰ��J������~�;�sF��+�G���/����&�jDdT�pZ,���!�:D�M�:Zk���ޘ����/�?kr� �K�y���B�&�R�7?�	�SUk����|����8>f�d�~�e�履�ڜ��Xː&<}�U�?�jf����K�_襥YGWjt�!���J�M=n!�*�3KIdde#�$a*����A��DVgK� $go��r#+FB�יr��!R�οr'�Y����:��s�	����p��g,��*��#Ne��҈<zܯc�T�_C��s�Q!��g���@J}�& �1�Ր��O�l_���ө2�ʫg��㺑mD�R=��#�*&�B`�p���Ў��?g�=6�X�.>t����%�w�e˒'�t����E��;|�c�çx���+��>ھ'�PLf͊�u k�VO����;��d���R��r[Ej����B�b��1n�|+�L)�&�q����Z���W�~���Tu��wH����ؘ?I��侁k1{���:��0b�a�讥v��S���z����]8 ��m�w칖v���Q��k]��^��oNO�o�n�8cD�ߢˍ��A�
/~��q�p�d�� 1>y��Ljh���|���x���I�uJ0ԶSk:�%]p���I-{�J�G��$-���G��k��7�| �@N�{�[*���d@'�C����q������Z��=�g�ҹK�{"z,�����|_�w��ڎ:S(���Ρ'��#��I_�x$7�H��ꖪ�)G�yd	F��tPì��� 7���Z}j;��/�]���ROc/�.�����)�� ����M�K�M�����>�~m$��YH��_�������/�ɕ �z�K$]ꫂ>}y"Ld�
�Dk���ךּ'Bc�?ď����o�qfbN��aK2LZ���E����ԭw1���.�J�>��Y�t�X+"�hEd>�z�}�u�p8�6��J��U�@�m��A� 3���?���������R�G������@�N��S��U�&�=���E�c{B*�Er�ӏ���	1�d>�x�֏w<8�ZG~�N�׍u� 0�2[,lB,��R�]�
���..�����F�- �Xu�h��]p�foXz�1ٛ��D�ϐc㎜kV�tTע�`��y�f������8|#�vخ@}��6�	����eK�.GMC��Їd�n|q[ގ�ֿU'���r�,SnQ30�.�^�^c�qH߆/V̽>#�o&*S�4�	9�42�m�)�x).L{� �=��4��VmW��4��4�5Ju�e7fa���&�	$�Py�q�{�����(����wȋ���<^x̲�{Y����L���"�ӵ�op��)خ.$���F(S$��bd~�y��M;umj;��ٶ(��"�RU�����э1c��\T��� F���w�����JU�N�Z�C0`��z�I)|)���a��V�;��7d=�六GZ1��:�G�ԥ�8SH�.|`�{��Z)۰GQ�<��}�1r�	e+ꜛV��|��O�f魞a>|m\w���K&�0��7j���k�;���8NBHb�TU�Ԃ�b@��0k��v�iǍ4�[>&4���=�΃�E=�T=j���$P��5A�])ݱ�F����@
c��-Xl; �T�DF�]���D�I���0k�#4�UN=�*~������)��('�@PUB#e�{8�#�V-Z�w~EH�MJ8��8��u�mmv5M�H2���&_k�M�2�H�Y̝�)�O�`Xy���/���cV���n�/�"6y�^�O�eC	���ޙ����2�ʾ�~/�/�������z�cc�UFp z�J)�Uo�H�����-;PX:����x�c�(��Fʇg(,��%_���E�	%k!DYc�t��t�!��̐���&�#������K(�D*�F�Z�6����[�2�>+�2��$�!
A��e	���"+��P����t}X����b���Q@�oئ�g�*�ŇF�eo8>-I2tXvujUL+"�R�c�T�LTE�����b4I����
����D���)��HO�)��Z]{���+c)�,q�Qn +[��(��	�Xe3ۦ3D�~Q��_�A���̺=<K���F���0o0�~n	��n/��V�q��7vBdE]�}��C_�@�!>�ܧ��o�k����_��_Y�E�6a}CŪw��G�2/¨��Ի������-O%��2�j|��H=��W����|څ�@���"���ͦIdB�*��2�� ���usoޥx ��R�����	��x��?�ww���?�*Ci7Љ�	�{s2���O)�G=�?���9^-��r�\�]�~�7A�`�K:9�7��"����]�˻�L*!�-i˷4,����0��^?���y��j��U���V����^@-��M����*���I�|q�Gl�;'g!��! ��YG�ҿ�C��x��\��:�`�,uu|!�p�pV�� ��^	��N�N�xD�D#�����Y������4+:���t|	Q�LbUGvV��BN�U�0���}�Nc��7Jd-QN��)��N@wrA3,��o�C9\��k����$����e�威W�0Z .��
7mP�����(&j]��#��f�P8�"������X$[M3mZl�3Շ�S��B��ڦT!&���ϕ"|�6�:~ͬJ��*n�Υ�0$��p=����u��,���BI�z�:(� �@pPk���[v9{� ��JRZ��V��Ƒ�1@����^��H��l=�bWc��V��rQٚ�O��C���^�K]�����y�w�?m�犫�e� x���"q��n�aJ5J�*[�*�[6����Յ��=*8J3��ᆳߴ@�(��_�����p���V�^O�:�*�������X����=�,Ҷ�n�-7pjc��7E_�����c~�)o|��H��:�b&w�S;��X�{-s�7*�<�ECx��٣��w�� ԃB����F���qn*�m� b¸��W92r~� ,+¥ȋgW,�ڍ����2C�n�qhu��y��pCP��h �����55�K�u��6���51	esx\ެWJ�@���NJF�`������)�/b_�e�@x����i�z�M`?�J-a����P� ��R,�ǅFK"!-����r�2�6V`�Z*z�f|N�g��e�k��]�9�����>�=�����	���v�T��=aH�o���(���R?��t�	�X7�x��L����CDE��s���R%�p�l�;6�Yu�1m}��%y���5��>����Z�k��6A������Y�v������-o���=?��7Sŵ|G�ar�fߛQ�����������C���H�O�%@b��o�v\�<����/��7a/��)d�ӓ��&�:G�ҹ	�}�芐0?��*�W�����J�:�q&��4�j�M{*՗;�&���;�-5���×Ԋl���_]Q���ѐTAA�?�N�=�9��tB�
��;Ѵ�?O�|u'�ƍ��CVY^!Q۫�[���̿2�wQ7�[l��W���b��y�E���?I��?�k@ì-��(��	�L���O+���VE߀�ņ2sc۪�+�	��ˋ�l�%�+L��Y���`��������O�Jb����p���%J��<���"�{���]��$�Cr�ΛQH���:W�$=�w�3���y��2eo�� ��eF/f�,&`Jj��zE�XM�]H���B������p� ���!7���Ɗ�&˴0\�Dݩ��+���ZVz�"����(_;sdT-�A*+���{��{y������)�<�K����W(�$HL�-A�+fiIFQ���B��{�H?�X�fSS#�KS��s�/�NzJe�������:ӱ4�
'qi�)x��g�P��zg����_P^��r"�C�+�1�4X��("Pۃi�GMM��d�Λ�8dA��  �G���R�ke��8�>���L�lҡ+�����%��pUsb�rs�))��\��i�
�*��o��y�{�c����a�y�bwn��Y�?�i��27H������S�BK�H@$~'g�,,� D��Q�<��w�Ȓ�B���fg�=�\�:����M��
�Pㄟ\[��e�^|!C��>���@yѸ������q�`��s�>�~�� !e��1�� �ȉӨI<e���*ZAj���1v�Hg5Vp c��,O<��I�H��3Oo�~�Tu;�����-�����Ѐ�,UWa=	V�����ɝ�5���n��}º2�������a��O�tY��,��|UJ��޳���m�����<��P�e ��K��K#Փ�'���O:�Jַە�l-§�#��ko6r"5-°s�UL�͊R#�t��2}���v�?�3�EnwࠤЬ�o�SX_��ފ��!T�p�eОꏞ�F�%5�����q��&8�۪�q�4�҃t�/���M-��,�H��]󏃱�?X� �8��. o�Ѡz��|DY�P,i�
Fm�K�D8���$�'�r�
�p3�c'�7�K���8�oYް�=i��^jh���Be'��Xr�l�3�i�6��u�0�O���W�Z�)�Y4g�O;�£~1����B���E��%_c��_bw�S��?B��`����5�z���#>����s���\D�k �We%��'�AI6�%�6kz���}�>�?K�vo7\�D���<��	v�S�5���7�F�|>������+��H�L^��"kA��|�;`��>��ߎEJ�d^���U1w2P�9蕜�9���K�6�g��Ozhj�!��@�]�(��D�		�Vu@#ȴ�7�ֈ\Q'�ʔ ��l��ça4ky�����+M�݉}�t��D���%
#�G�ر��K+okE����B��ϨU��d����A#ӝT�L��t͹���n��Y}��
��KW_ �0�f�2A�
`[H~o��IQ�x8�!K�Տ���]�35�L�oah��`6`p���Gj��+G{P\+�M0�%e)�ī�`�G1iIaNiI0�^�'��c�������Y<s�	]�H�/��~���JAĳ,S.�W���ѣn��	��M{�q�\ڋ^Q�ʗ��Aݻ��@ En
-�a�8R(�M�"3�D�`�ҩl���t��+MU�5$��X�nz����9zKCͮ��lF�@���}�}�k:�#\>̔q]��e�㭢8��!o�W �/X9�XS�q!|��=:��A��Y;r��y�^�խ��3����=�š�)
�"��A�X̺��ڳ�k����Hl�Oý���z����^��bu�a��`s��;Ag��o��,�Pl��2"4]Ы�����Hm��Q�{��~�:ص���c���Q��&��d��de�y��
��2|��DL��D�#�u3��Tʄ/'�$���"
A���A�B��S{re�OZ!޿�8@>�3�a#V��O۰�C��������U�6g�n���@�v�3���N�\ڤ_�,ہwE7���%Lc�W�{�寂�����q�e4���ZJ��F�$w<���ay:��Фc1���R��f��m�4MK̰WPAh$�{�������Pа�±���=�F����ˉ������)荲���8����#y3���"��[�H,�E��ˠ�w��td��R(Q	Aʓd]���Lx$��͋�C�Mf=��'�T�O9^ػ����KP(����
�B�q��Y�[���������Ͼ�v� ����~4c�����,d��
ɍ����Z2|9��+�2�f9�=��6
X�D�/l�ķM�7�q��)B��R�t��:E������}a�b�}�0�Kt�D�ecgv�� �x��v�C��hB�!���}���u32�$*
�kg�2*8�K�����W�kx��P��6I{�?���ᶂpو�l�N4_I�gRo�%����W��<�~����*Xl�[]���մ�L��N��!�wd�k�,K�;jk�{+�`׫	��o�n��ê2>���_6�	���G�}c'	�������.��ٔf���G�m�hDvr? ��e�����C1~ϒ"鄮�?�S���#x\y�Ҳ���I�������Ԭ��I$=l���$��8X���	�.����^��~�rify�5����V����9�إ�޸��[�O���*�8�ʁ ��M���A7Ye�:�ഊD���(�^�?)Y=�|��U��}ق��Hg[gbU��I�%�OK��-�̉\�Q��|�@�;Mʙ�V��)���#w���sY�I<o��0���(���0+Z�����R˽')%^��qb��r�[�[�3RyNsяH��E�x���3���K�B�lJ�{Ӌ��v�NW�qŖ]h��Ye]@��9{;�By3�Fxh�W7�s/�i��J�I��d_e���]�~ij=d�����:�=p�8�9"KBEtºw̑i���.�A��[��I�b�5��z�|Z2��ɧc��8r���&n/g��x�T"ɹ78@d?��C5��R����/%L���ַIo1MF�%�c,�cb���Sp��<%h������zyç~����1I�k���L�,����i�#�W����uꨪg:�Ȅ�ޔ�����ê]�,�����%�u�:DA��#����2J�г%H2�����wǠ�������J@r5�a�����:h\���-�.��BCߚni��ϙm`���D�dɏƝ�/��R��tk�� [|���+��~D�4q<���|_8;%Y��eX�飩P'�V�VJ�m��!�jTs�%�	���>�M��_FrqK��D��7�q�@�f��g)=Ļ��sɤ�z�S�0T-��Hw˯�H.���q�YO����<"���sR��Gv��b%��Y�j`��F��HV-��z��̓_���������mo����kq���j��-�&��M��z(Gӊ�U�(����T{_���!��2��m������	�N����`o�S^YjgmܾT�vb�7�D�5.��6f=�ثS��v:݂W�#����꠳���`��dmU��FO�z�ᑨ�L�?�~=X�d�_���,e�k u��@��k�����x]l�.W�D���7�i�T��
��72�� i7�VC�~y�z��;2�����-nS�ޛ�\�2�C+ iT�����51����6���rw17􄑇�&JFA��[�W�3	D7�<J5o�T����C���sTv�����aؖX��h8���q\�ԧ�,A�_�^��ɸ�A��Tkg��cF�<P��$��.]�-��m � D��DܙN�8ǐ:䧞�=�����B���Z肕�{��B �M�(��5��\:A�{�_S�~��4C�q:"�qוH$Y�.b�A>���f[���.j�/���JO a����+v�~���aM[/��u��e�N�B{��#�8T�N��}�B.ч����v�)���o���F���T��4S%��������;����f��q`�&t�A�e���(ϟg�]��t�l5C�����HJ���N��*Bbu�X�j�n�y^�?f �imoQHȄ�%����q�݊��A1��<J-���I���$�	V��P�ݎ�:��y�L:�LEo'���G�T�D�܂���:�G5��Y�v�ŝh�T{/���P�e�X <�4]��ۥ����-�UB�j�&���ڬ�z!��LJ\�K"�N�#��G��d�%�.�ުQ~����p�"4�U,3�!��֌���������v4�'�c
�����Yc� �>�3�B��#��4 �+� ��L�����q�K��h֐�8�����~�ʉS�Y׷h��T��
f�n�<�X��B�.l*��77�oٟ�iq3��)z�~��zM�*V�N������e�6it���aaO��&�0�v��P%�|�W�ď8����T�3Gr���
��UN[���Mw��#���?�Dl�)'�I��2Ӧ��]_��E9��B'�M�kp����R�B�w<Y��n�MJ�u�"�Xz�Y�iț�"��ω�h.��W�z�:K�.�Яc���,�Âڼ���k�� ��c�_��A���rL���+�K�h�Ew)\��#�Y��D�,�PO4T�!c/�*�i���U�=y����i-A���[d
��Rq�h�n:�'F����l�s�-S4E���kf/��g���e���	a���!o0ڑrˉ���ĜC4��I�_>d)|�x%`&��Mj�Ȗ�����]�O����U��n�L�3��׊@�{BZ��Lt���GC��Nw�y��kY�wn%����f��ܡ������x%K���Q䜉���+��"���?R_b*�2�c(Z��u��A5b{f�V*/�*�.�ݣ[{��率Ή����v^4�$E�L�l7�)	O��"�۴$�:��I�Z��F#�L����āGh��<�Rn׭q�!�׮�"\M��� Qݧ[�����j���_艸b����(f����!�%�a޶�y����C@A�ڃ�~�s�` [�`�"���^�%p�+�PAM{��ZY$(1,�th�x�����0��_b�/?��J�)����(i������U��xQ$�en`�sN�b
,���P"w|ǃ�2 ��EM����U5B�D�ddat�e�qJ=Ȧ��2�j��+��_�Oul�h*��̰�$����xAeX�sQD=~�ƚ$ ���ܲJ�Qji�����ҡ�x�C[��H\PV@X�/�`qc}��^=���'�m�~?M)B�����X���.��)0��d�j]߬9�eO����� H�-6���79[��-�!��d��Ze/iO[Ry����!��T ?�-*U�Y6}Z�֡3�x�2�'���ꁵ\O��`�����3Tqm��L� (���nE ߓ� EA�7̱��>�-�q��6{�Mh4���U�*j�BļCQo�P�8��ۯ�Y����:�3IN�wِf�`��ʿ�oN��U9��C�l+�]i�H?A�D�S��d� �޸T|XX�_+ZD���f�/G7�c���.\Ng1}���%�A��t��0ڂ9� �唒?� �i2'�6�+�O ύ�x�+�,1ڸ���M*�a��V������u�O^[=���b(�d�ζ�#�>Ck~ÛQ�|�q��U�b7��Nc��{L�	mݸ��N�!�i�Uj}�[�m�|h������Mg�ƪ���0 � �����o�H	>��K5��!�֯�C�� <4�A*����[�9 rƵ��{pQ�g"�Ȓ�
Fp4���B�ʊ^�Q��#�9�1	��FR16��ײzmP	=U+���)��x�꣛�?�� ���简E/�ln��R�X�vg��_���������[��_�&�{�ؔ���	R������
w8m�:�D	���8�~ќ[�CrFT���$�����(d�u�E���L���&
����[I�]���Ժ�f�޻@Bs�6g�����0�q�5�'bs��o(�$��k��tJ�4a$�6K��zW�"�X�N���'������oA�h�Z��K�%��8��(�ϱ�"-n9bJ;F���Di���kY촦l5�8L�FIw;i�ఱ��:������d�ׇG�� ���Ȯ놱����f��29��bi���s��
���<5�''Ӟ<(�#���y�?��p����%��X1�up@��$�S���َ&�,?t�9j�*�޹l�$���G�b5�j��Z`��i�il��r-�e /�<���y.����[/����a����/�b���rk/�6@V@j�)�yUy��|��~TC#5�Cx�
��eC�}�����g��ғ��:��hUh�p����RO+�_�)���[,&ީ��u�\"���vl.�K4	���/^�'=�y�L��������O�7 �?g�?�$���{�� �B��?�OD��W����F��t�(Ե�u�]�{Q�D���d,��FȻ�������q12�)�C��.g+Y�84l�K��j�E��
}s�9p\�p˒�󨚃|Ȕ�u9��m�_�20�}ͮI9o�7ehס�Qb8n�Q�3�暈����#4ӗvA���o��k������K,��ΐg�D}3x+-e���ߌ�Zm���9D]Fe�nitE�N����1�8��������Q����������M�S�A3hp�O�J$�"3�Fo<%|q�z�Gƛ[烜D]|��fH���/u��'�7��?�*H6r�Ht�� ���8]�����.%�">���9iZ-C����ꆍF��.X���
�T��V��J�gE|����]+O�)�/�s��_�B�dS
6�혣�C#r�ܻ�W�A`���M���ݵ���Hte,�������*.�O�b������'2��k��^k~�Vx���'���7��fQ�+��wР'���P�ATf"�}�Hz$	Ar�{}#?�v�"8�Կ�P�"t?��]暗I94�x���M�E��m�����壋D�1y����|�Zv&��k& ����!���
+es�v�cU*c_�8�@���N�Y<�R,��s� ��o�qsp% �6�]~Uu�ut9����N��$�]��-�����l�X6��W"��d��Q����ي�4� �j�45?jDڎ}���E�VlK2���c�����"7�L�k�A�D��'��l6���B�B x!�Z�F.&nj.���d�܃mt�B�I�[9?)���������T�.�k�k��<�뒹�(��Q`��إf�I���i��<��;$��N���{-6u{V�S�n]6��d[0�V��cC���SO�]%P�2�(&��aj���]¨�_�@��n*�!�`��7�
d\>S��M!����y�V���
��{
��r�JQ��� �Epm{"�gLς��A��Ea�@�ۻ"t��W4���\��� <��\�)Z�hʳJ�3�^N_<�[Se垸�^����!'�6NB��������W��d5�D���-w�
�h��m��Ӗo�\�ɔ�#r���&�=>`�T�c���+;�p5�O|/x0��E�X�y���&R)z��itq�x9���Ag�:2�[ ����ǻ�짒�Y��? �yP��&�I}��X�<l.i����M_� �]�u���SB/3㸚^['zp��P�B�hL�[,�W�/�=�֤��/n�0к���n�m����\rd�Idx4�םf���SyA�@�,�v�d� ���ٗ,�������`G����h��^�@�ڞ��8�*6ܧ�M���Ɣ�/���S�Q���(�)��HTƗRoiq�%D���F$��64��t)�y0��>,�]D>�&���Z*�:׸���`��>Yܕ�z-b�D���	r�=�C�	B/���%�`FVΘY�]�A�s���B��qȐ�]Yi����t�$L����M��X������Զ��F���L�t1u��-��M=7*��	Ȯ���zr�~C���{Ѵ1c���~�:�/��&���"k*���F0�B��;��b��-:9��[zF˵���d���xD���L�[%!����,^ҝ�^�y�Oo��?��|0��ٷ�<H����� ��;ǡ�B��n�Ϝ:��JA���. �$����Y[?�H�c4��j.�V�$l�̹����z�c��2_�"S�0�N�7i"�ho��q�cW��H����^>J��K���m������:�>)d��QY��6\Q�d��)7��mT��Kg�*���T�k��(�}'_�W���h݌��� c����a7�rZ��F�D=�Ѕ��e+��ڗ�x��� �;ևQ3�(��bS2C�68Rs-�X��%<Us�Ԝ��³����~��*�-%������d��B������Ə���v�c
�w@\}����ܗ����8��~ɤ�)o�uCj�J�,>x2�"[�xl�O+H��L��D5�K�y�\TM�W�w����|�����+nΗ��V+�J{�$؂12�+���������D`n��3H�HY���CDf0���{3��:��N	,�!�h>��mT��4*�@҂������\�&�99]�tN�D�]	��°������Gn�qEH=��U�w�*b�Lc6����%��9�8������J6���!X��q�y��~��ڲ�@�GF	hp�]<�rd��U�w���[��^��|܏L�"Bc��z*�W9����T�V�ZX�f�x66�������%aB{j8k�H�J�`�������_�5�خ�Ę�`��Ʊ��UB��!әQؙ���ٶ0�����s����Q�X������R�A�V"[w�^D>/Ů�:rmu�ġ��.�Y�3�?����JZ^��<_�tp�7gv	���Ϙ��� ��q��x����JQQm�EJE#��K����^��!���_0��W�[�4x��f�e�US�n~�o.ruU��S5���-��6�3�8��%��/�������t���v�u����;�FA�8$9��v����Ikw�!�T�
땀��i��v9�x ��y܊u����yG�����k�.�ſ`0��O]��-|Ɓ�,���*����`Ï�W&��"B<��b�3֜l��f֞ų����z|�g7}C�o�\s�f�?��{���B�|�ni�>���>�Q���ϼ������BK�Q�R��������_+[�4��D�������b�џn�ꆇ�Y�C�SFO��SW4��p3���7�HL6*Nn�q/���\��Xpl����,H�> ��1��N��\�\���!�i����Y�C�o�����w	pD`����a�ǆJR������.�,�k���x�*YW�NzDA4#�{�D��j��'7�����*avo�(�rs���~Y�4�hܖ�
�ug*�1�rgQs�(��܍9�X]�|ax��u�L�M���I��Np�
!e����a�ܿ�Oǧ���.�
XmA���+f�"��lfS����=e%^<��n��pD�F��kB������'�5w��^�<pM{�Y��$)����I,g@P�����h
�hK���>� cɯ�x�i���B?Ʃ7��M�B�r��%w� '�����߀o�[���\��<��$�vZL���Fv���d�X���R�UB�'���@�J��TpqvV,Y�d>��iw���O����O�[��jѨ�r,�Fh2n�o�m��������v��C�Y��i��SB���:������d��q2�%�+��q�YJ�2Mp���K��#�H�N�'�Q�&��k�[]C��N�3} �n�$:d`������m��\�P�/C�{
;7�n?]t�+�{��@�����*�� �F0�T�D�a�!����(� ��	rȞ|���S�Nڕn0�*GЋ̺��@Y�AcqUŚ�)w��5�� �;Ά!6�#A1��-@&35o�W��z�D��R�N?���@�p����@�ö]bvZ 	�4��Ӊ4[m��{^g{�kX�E`å� g ��X�e�������ƖB��*��m+�.����DbY�o��J�� ���� (b�.��|� C�_D���*�^;�k�C�w+83 �G�(������܏l:|6vnUh��i���·*�o-qív�I��c��=�;�����^1@*�
���ѳk��$`Rx�0~�.�';�������M�tt����"���	��J���X3��d|�6��K��#u����M�7]W��ɚ��Z�e�<K&�푪���'B���ͼ�.��ST�M��;����B֗dԘ1����tE��n_ֺͦPn��FR���H��ozz�X,:v��{ͩ@�V}�����X1��bZ�f�6��ZV�-1���)�@q��Kwl8%)�!v�ܺ����H������O��%��Nx�(� ���Ϟn���Ք�?U*�ÄX�1iX�X�䲣���I^lH�ub=��Ҋ �rdr4��=	~�n�6b��<K�t��ly� PGҕ��Q�2<�g��:�Y�+EXi�fP�������sV�`�6Ĥ�{���XG�B�����_ZAe(5����K��������};�q��q�WU������@�\�*W�m.���w\h�Ǖ��<�MuR�)�1I��z�#����=�d�Y%9l�t�
�1O�����U�1�T�'FnIecx�H��6=mE�{B>L;�2�&	�c�kf�$IV���������ml��(O��yn�����Z��i�u	Da~[xk�W�O_�kA��ەE�J��Ҕ�:�x֑�TżZj3�:���[<�����|NY�_�Wט?���6���FGY!L�,~I�a{����V�{��R� 5	�����ɉɝ�<�R���Ig=?zI:��ү�r]
 ���\�;o5S0�n��l$��]ܖ੠D��V����G
��m��M�3U�����w6�W�2c@ǍJ��b�q�V���Rֵ��e^�b6�\u(yo�^<�T`��l�����v��'��>-�4��!Ò����N��*ʕ���0������(Fk!�[����)ʅ}�@�N�Ҫ��ʃ<L�H�5�CP���a4���kH��Z�e����6���q��e���t'7i�I#8^v�e��F�UD�CU�+����������N9�b�⪪j�S���T���� �YRH�u�;Op���z��+����-�=x�����__�V��X���:�� F��r}.y�ms�5�؇�R�(�cq��O�|����7��X��v��� �m�?��g2��Ʀ�%�!��1���&�:3z��$�]Z�f�$���7<��Sx���;�}�`o�F��*�������lvF�8�(�����tr���)�������W	�D0aZp�Z�ؤ(h�`�/8| ����¯�ض�sYY�i�s�����+�j]�
$���8;�iU�'�{����ռ~��Ch2g��C.�dI��I�7�J��z��B�q�ټg!Z�eޟ�]�Ib��j�27�BrKC#,��hd�T���q��Q$��My�2-2&�0(�is�� 
�N���7�M��/��Q�AI7,�g�Ag��M I1�5N��瑗����*�m�X�!wr�_��^��IX?|�TA��	{��<�j[,��m���f�0�¬\�^���t�~�P��-�N3㠇���
bY,�l����+8y����=c����=cÃ{Bf���4���Z�C�N���o9E�m��k,��Iq���u��h!/�e�z�U�$�)�x�}c������?o]�t��8)``R�|g��Pq�s������R�1��ޱ�+4��']Q�"�N���7x� î=_�2{ї�`�����q����!v&;��hF�F
j�N�%�(F?�;�|�i�l-ٻ0|���uyC����������
�$ +DD��˛� ��!s����\��2��q�Ew�g���xA ���Q9)a�&w�E7��>���8\']��R���k���{:�A�1Ƃ)�B��ܲ���S텮b�J����тɼ(i��մu��25^k��������'&{���)Q��|�iM���A�:2hx�ҁ�ܪS��<�&mC�+NlqZz�2H.�b�b'_]��Nbf�� �����hf�qlS���;^5�4v��s�[`����9���xJGMg��J���:�Z�[8���Pg �V[]�g��� ��3��O���GTl�]b�C҂OV��Xef/p�%�b�_DtM��C��
*���c����w��)%JҐv=U�99-lpY(�E�/&���}ΐ�,����H~��A��cWAZިX�Q�q;;3g�٧E�����'��D�j����ؕ-��O_��s��`�7�u�>/kқO�Ԁ�������·�����#���:�a+�����z�	,��FZ{�+�77'�-��{�u�mr��Z&TI+��e�>�-.�N�Y���D�uA���Z���&/��/��$�vU��gɿ�!&	jTk��T?����$I߇wl�����p�z!�|\��آ#f�-	��8� �I-�`�o#=��S���q�RF�ƕ��J>H�:�W^C�[P��? #S�E�Z6��ʗ*�Y��o�[�/��Q�ĮT��9�nw���?��,���~$mO=�'[w�@�ZL�>�f΀��~ 1�������y��`S�
n5���U�s���ܥ�~��t�
1ȃclv��2쭅����0U����/���Rn����;t�?(���ǀ�3���h,�}�B�y;���#F� ���Ծ T���F�vE����&]��_S�(C.�+��*Ih�~�E��߼�'N��y(�XE�����Sޫ�<�������ہ7���]SV�r�x�����JPә�͈�(4齮5���o��v�����r���ay}6�P�� �@�qO������6�b�����2"��D�O��8dj�p_BWWa������/Y��=D����M(
��-p���܎����?1�E;�V"��ą�4z�Vg�}��Ff�X���z�M{z�P/ߵ,P� ���k(�R��P)�"���P3y��_G".�lX����SݬaHL�,�F2M"I�p���<}���H$휝�+�!�d��)n�S�m�%[t��GC�nA�z���!X�M}{A��޺-�����nE�:�H����
@[쮋r�FS1o5�
��<r:"���%Mwna�U�Vc!M������Zڰ��oMͥ��L��p&�aZ�1hĒ��'�n��Q7���Yw9����e��0昂�ҍt|U#��;�ɊC�P�W�/��Б_�+6j�lQ�ӅQ8&���r����y�?�#�1�&�j�:��Ca��`
& d��"9,�b�'	Ͽ��zW$�$+OIß��-�ɵ3�y��Y�.�&vEq��
@c]��`�%cȓB*!?�3���B���e4��mK�m���*f�a=]{�MTNǂw��r���Y�� r\)���\?X��1���ش�^@~2�ʿ3�|:���fJK����6t�Q5�K��E=��Z���nT��^��#�ڡ�t��������i=Hu�0$�J߻�vv�X��u�"�a+U��yU�h�����{I��Q����v��ny� ���t�o�I�ǢHW��U��C���%�zs��}�n�.�w�k�a�1ם��^��așv�c����{�>@`M�T���O�u߁�)��g
Ym�GA�g���͎:�����~m�pBk�m�:�����)��`ʐ�mS��(�\����=Q�$�h2K����kƾz�t5��D�t�7f�d�Xu/�^K-��J2Q%n�fw:�D�ƶ�
{y�Ԭcq*X�ne�t�/V�+�^��7U���+��o,��p�)����2
��JsAA,�a���s��e��WN�[ܞꙔ$�'�#��n~�$B���C��(^��ẩ��i�?����c�g���k��Vs$l�(3mNٻh��J�m\5.�jB3N��1��c�8q	�zAYVy2��JB������5� ��Y`z7�7p��s�AG	j����_��ƞ��a��yDoB��V�5�&u��.�k�0'B�?��4��@�F���e24�-�;\���~��F����T��˞0>���`%�����h����#�\�	��&�5�Ñ�VBykۉ� ��������e%�̔���j`uZk��xTud�PPT�$$G�`8=�\�S|���*s�ل������<j���׋7�λMf7� <����D�����q2d�̶�.�p�,����ח���P��\v�JOԶ��J9����F�����v`����2M�eKi���1t(��[��o��F��	P��ͽ����+ݢ��eZլ����c�M�;�'ٰ���<���Պ��4E�o)^ԛ.��Xȣ�?�[X�X�1�U�
�J��_w��b"���i�Nͬ߈aR7�����	���*��!���e�Gc����Ovz�rCA�0�sa�m|��OL�>��q���W5�V���N�2���lz ۪�=/SWY�~!��4�L��Ն�s]Y1��I����\��= �Q���5ڜv-��V+��8�SLT��Q~�v�B5(�e��ps���Մ@��$���n��bmGb5fD�~����/R�UIn�pH\��`X����E��/T�J��T��:dO�^���~ �R0;(^]!�{x�^eތk�ow�ݎ�ɒa>{�:k!p3RdZ*Mjaq�;!�!n�׌����VW�0;'j��X-���r"��s�r�vf�0|T��7��E�f~�t���Q�ޢ2z}XU�&-PV��u}�h�#��d��J+9�t�� Kڮ:��~Uz�<#�4g��9�6�'�Z{ &=3��y_�ݕ�������n�'�x��7�� �*~�D����c��IH��� l�2n=ai��$Y'\R�s��Pm�ۥj�2m�Q]�O5�p����@�o0��'��<���tP�;ll}�����^�T�]R��6�^��.BFP̙���f�"4�h�n%�6 ��3BK���<dˏ�B#��}�v�O��n��@�2фUT���q�;Z��Xx��� 㾄 !�f>8���G��o�*�g_��	��ߍ��|���^O�G�1���Ā7�Qr*��BI���N�d��H��T{�����\�%�K@
�	��s��ݺܔ)AH����c[@MǙ=%+� \%���vD�tK�9>����HR�I���te��Q�`��!�-���h@�X�k�.K~�i�d}(VEt#Tv1g�7؏r,��h����������޸:��}�{�%I0zJw����������c�o�����KE�ٹ]y��$�	��ngT�dmR�Bg�A�e-=Л ��T��Ca�Ӯ�{A��]�up���af��s�<���LIl� �[�(Xt��J�0P�	���JC8�i��q���o�5��h�l�}�!Jr�,�+�H�X�ܮ"2��"�W�F�~��������s)�=���Ǜ���H��*$�.�n������>�'(����9�?��p�G�ʾ��C�
]��m ����Y_lk+��v���~�8�ϭ��um��f��̍F�^%��VOZB��O�J�d6���?�����vm������C�(�����s�Gg�D:���,�$`7�)Zװ5�c��)aײ�t���J߹Z�m���TR0�Q�R���W�՗\(}��e�r����q^��YNW��7L(�>������1�df���Y"[����.�����)��0�d(��� e|�D�������fϛ5������B��q�䊉��T;��`@g�cWB����$�
�	Ɏ�KKX��`b�`��B[ '%�����i�=���{#������� �p5}�$s�$��d;S�Nz ��/����6۰`1�v0�h�˙WF�A�<`�r�9�k﮴�.]=v_��~�TbIj���D��s:$+^Θ�["��Ǚ/������2n��$��ó-ݳ}$Wʯm�u|�a�K���=���~[%2����^m)�ԈxU�j?r��yi�3u�Ȱ��s
��/EW�"9�-�l�gw��u�$�}H%�}�B�f}����Ur�\<�g(��6��/2x�(�E(�^�h��.��*�`s3qJ�!T3��[Y�!��,Em�,�c<`�c�x�����r�_�dtΟ���C>��p
Q�B�C��)t�-ǭ�Z����F��W�ږ1��_.F}�t:բxသ��[�V��?�@�3n(iS��X��P�f���ux;
���5(�E�:b�1L�x�[W�b�v���
�W�L����f�u5$P�"R$�q�{����shN�(yc��� ����1G><)�rZ�O9�0�'{��q�r�D����G���c���[T��岹CY��x��*�����P����M"x���_+����|ϻ�(3���$���ё����V��}�m��1����52kY�>3��W⼟�n���o�o����W�l�.J�(�2tx��#��!9�S�WIVk�� ��e�T����S���26�ė{��!���������p^���S�R}ʽ�S�8hq����}14z�����6��G��L#(��\�����{a%���!��1���_;�}ΊNb5� !l�HuK��籾�� �������%P��������u}�4K�8C�s�&���Z�GL�����-�S����Zꎻ^�H	f�^�a�#�E���*V���لG3��Z��t�s�ĪT�m�����xj��YP��W�
�5X��U�bW��	S�xW�j3C�|Y?C��e~W #�\^m����=3E�ƣ6��{\/����Ί����xa��6�u_�@7��3��f���R�!v	*��l��a�<��RR>ZmE�:o�+��ſ)�L�����v,��8�)��"��@rh�� �?ׄ���\�C��p>D���Z���Wyx�ƙ�:&־�;A�b��d:Pؽ�"x�|=�O��E���ѭ��8aU�x]U�%��ׂ�����5nv.M$"�[�aB��B�x�*AO�5�����b�E6F�ȕQ=�f�C.늹� ��1�<�������uG�3�\� &L�q㯁�V� �b�>Z�~Z��Y<9w��UH��7	qS���{�|�<0������8�D[��Z�"l^��܏�&#Z�ݨ��P����(�S��.������,���g	��>�	A-&�^%��8�EnQĲ�@}����x�����c��e�1ձ�n,VQ���j����!Lkr"���ݯ�����l/T��;�����5ƚڛ�r$�.H��p��#�x������\lG���"��f�2���ԫ���GSĂ�ޏ��Xh�L���h�ٴ�MS�Z�i�tcNKQ�g��q���d�	�r��˞7��b��\$�;tQQ�\��w��dt6�^�<��Ex�Y��f!0�/��h�!j�zsd�p�j#JY��<���o�qH��IP���� 0�{��Q~�<�gt��l{���~0���$}U^�_�v����?�q��ST5:���`�D���-}Wv�q����+���2����������(,�x�� ߯�;��	晸�$,�)4S3�6E[��wp�b��?dȠv�y���Q!)(�.��iPr6�u�����Zxs�IBʥdG�����.p8q0}hy=�z�����6m������P��Q�R��E��2��V'�@�����W����	�<"��\?(�A�Z|���bv�B���m�Ng��8�[���O$�����b3Eƭ�	橖���Y]���?VN2",aรC7$�jCw�z���>�*]l0o`GUI�=�%��{	\���/��Y�2���XB�W&Q�MO��ù�d��]��
J1�݁,��e�m���,�Œ�X��կ�͐�F��(�����%�?�e{�Y��e�����K�)�A���"<:���=�p��K�M�}oτ��h6xCRnRWb��E_�����'�%�M�}$�uP̈́Rpez1�����"�����h{��5$̶:��M�6?�3#B(��c�4�<wu�Nn|@c��Au998ԡ�<��Ec�~M�W��*�T�m�N�nc�Ì�Y�-�LLنH�!���3P;i�"���T$<.I�.�b�UIv���~W�����~X$�)���<Up���mͲ2vf�S?�����:�v�쮜Z^�5�<�S��9�~�dZ@hÞ�j�Y��[��-�����+�7N��x8�9wKuvB�}��'.]ūG����s7�R�qkKU��0mKV�?���6��y�B'���Fw�2u_ڏ�K�������űTM>�a��]�P��t�X 1pbY8M�vN�~Z�H�ω�vV�՟i�Q����Tv�j��r�I� O���}��,N��ɠ�����G7�tO9���C������ø���i��B��~�k;�s�����ٵK�ϦTJ�m�`���|���dr��Kn�Qp��7�u�h���ګ����B>T�	.e{0,�0�~�����5��#�t�[Ev0)t��X/
n�b�J2��ve+�Z�'��bK�g�Z:R1�mKiR$����%Tifʆ�
��Ky�
]�x��u:���
5�Ɨ�[�N\���la�PQx~j�p[̈D_�|J����(��6�����;�������)l¨\����HE�4|}�3:��_3��t]�!�v� r�M�e���6�9ǑI�V����:]��̀S�\$�j�{��ws1XK��i6XN���;ͲL�ɰ0��[��&o)�Zھ?zu�yĺ��L�%x�Fn�,��?2|��&o�kS�#�&{K��
ʺJkI��z�u�,��J��0�p�3�+d��pU}����kVP��-K�6!c4�����lBӭ��d.@��ƑZ;ʹ��l? jN�+c
���/��$U�^����[�߲��>s}��Rg�V�jhQ�M���!ekm�$z)�ȋD��!VX���T�[=<��jꏧ��Ρ���H���O�í*���V?���s���KX=̊Mq�Ù�<�)A�&��n5J���%�0�|�E-%2H�B��� �$�j�^�tқh����:��^�eD�j{;����9g��hZ���L�{:1>����dD�̀3�]�}~&�ɂ�^̃����g+D)�����|qi���r�N�]Z��$�������qr9��!�`��Y��&׮�t�e���oF�	lV?%!���W��n:�Q�����q����>]@�U� G��3ɕ���e'�z��(�:Wn.�Q9��GdQuR����T���4SZ�wf�;�d�`��^�	��5��F���N�%є��X�,,�j�T|zpk�Nt,�G[�,eLbQ�6X��{�)&D�}�=!�P�6w1%G�#h���ݑp��$M����?�u�(�H8�m�r��Y��StY�����N�v�ɀ(kL����H��u��L���y)`�?���B[J)����Ӟ��0�!� dJ1�Mb��4nN���0�2Yh��$���=G���6��*I	p+���e�MQ�ݭۅ�>_�I�	<����)���e�yN�\Z�H'�Պ�2Ѷ��V�JT߃�^&x�%���>����[;æ@Z�^�=S��0h�&S�)%�0���贇���)� y`���e���P�;w�]�~�&�mù�q�����+�4�7�����W����e���^Y<C�"�D���w�=�*#�6����:,4l������U\<h�\K�����Q[0?(p�~���.�e���?x�����X��6��L�����^&D��\KN@���O[w&H+�>��{l���Hs�L��q��5�s�"��針���%����WI�`j�l����}P�z�6���g�ntڮ������iM��������0��}
�5��L[�fb�{g H�|��&�y�j�S�m��Y�$�b��<{n�彤ݫ�+J&�36��3�S�jۄ𑛻�[�N�%����x���T�ÇG��S���,+UY���4�A�
�RU��jx}�S[0��V7BXF�13 �|$��M���H\u�!�b��[��,\���d��-j��8c1+7�]+�z6e����C%���|�Am˘�s6U}F��!�7+wx���_�g���b��1�)|��J����M�v�(W�%t��^��߀���C�̄s�; ��Uu�c�N>�YJ�C�0�{L�,���<�#;���ݪ���FxQ�<��48�ۻd���]\�β���! �md�4ܻC`��Z�B�_�d�94� G�S&%.�CHE3$�s�P�O&|ɿU�"�T�8Mr~��!	X��,�u�D�2�R���/�s����%D�wĒݳd�M������' �F�㗲c�Iu�d!���mf�>&���{=Y���ܪ������  <�?�s��#\��W�	�Q�<�ߕ��N�c�G��������j�p"�F?F[*� n�`���"(9x�h�>�o��5ŔF0%����ԦW���D�2�ɸZ��"�@>r�C��>"|��0��	G�d~.��9�ZE�}31�j(~?N�*=|+*D����k8�/���s���+gN�R�Wk�-`Z^_dڬ��HF��pƵ�I�����\}{D6D��O�誜5V��;X�B�pl6��I�잘\\�"	�W ��si/^��?In����^���>O��W!h�/�Mլ�T猹5�J�^�;Ics�<���ZD,�A�0�3�����S�`���ֺ��0�e�:�� Z�p��+�~SΕ���[��6��4f�<�G���8�4�@�Lj���i�qeB?&���עґ�5���5t�1�����_�N߫�&|x�[��G6@�Z�s$��5
�Kw�@�U����V���W���?o� �NbE���8A�z�a-� {D�^���h/.Q�c�V�������J&���Lb�XܥqEV�uM�i�n�R��o��t`��=|���.�)f_{�U]�joIL7�tj,�3V�����8��hإO)����]�0��Ib�/�i�O�G
����b�an�m� D�^4g��/��9"�+�"D��[V��]Ȍ:��7�*�����aP��d�}�6�q�8�@����U�#�����AO�[��$��񸙹ǩ�{$���ط�8���[�#>�h�	h۱d=���j��M�4��a�g���PfY$tw<@�7GwsX6�lԢ0���P�nϝ#T�F-#{@����'gKj(-'w�(�</�����`� ����n�+c���PT=;���D�����,5���_/��a���5�}�u�7����J�:�g��xH~��B��,	�䉑$����$�p��o�t�*<��HT;:�@L|�)��؈ "�!+�T�WK�����Is���ǅv�y�/5�9<�-�W_�^��8���N�?0F�1"�"((2)�$Nr��Ru8�I@��_�e�[�v�R̘)T�tuK�!�ty�7s��JO�Fn����5���n�!��A/����oj@[M�_����K��K��ڗ^ť$�����z��e��O}+S��oD��O�C�ã�sY�
%L�G����(�ސQd��U橡�g	�*�ag,����������p�O͌#'�ï������\��A�R�ᇛ�X}e!�N)؏�x�;K�GG��[]RSC�R��^��1:�	�I\�����?�E���خvr&1X6\VIu;e�R��_oN��s97*�zG&�~V����)չ�/=C��c�x����ES��c�r���gC�!����a���5�B�̐Ƒ�I/�I6����5	v�W��a�r��Rʟ;�����\���jyG$��(�"{�v�u�
j���O�LT+h]������hG��=Ksţ�6*ج�Z�������n��N����.M4�?��r��ׅO��U($�����a�m�}dv����63��8��m[��¬�!��U�6F��h�Af�Gpܕ�a�S>�F�<��Q�|�K�0i�S]������<���s��D���5�vl	���(���i4Z}������,.�;���;��b����?�;�mx�Sg<b䨩/���yڭ���w�6᧘N�#�C��%̛$��1�с�_c�1@����j�&
\����#�����M;�����2�S��Kr���n����ϥI�C�T��;��(�� �xt7e��.%� �F�jw�զ0b_�bإ6H��M�5��Y�o�$��(^�
� �� G/^q|cJ��'T>�Jj�0�L��Ậ���w�`ٶ:>�䷠��I�{LI:(K�'�
����IO�(����H�r��n�P���������S����D��FM���iV$��m5O�Υ;(�Ӥ�7;+Y�nu� �T*%"��)&��6Y"/�D+C>@��� ͜���d{ԍ�l��;�lN�����*un`�n]I�4/�oڿJ"1<��1�0s ?�T�#�<�cٍakYg�j(LB��m?󦬦AKOVY�P����ff|ڭD�K�JS&�;7U;��5��>e�ȧ����}xe���oXnO^��瘯 �9n�LDFP|�K���ns!zki3��pR��IJWG�m�t�@d`��,K>bKL*r�����������еM�S�v���{��_��G�l��$'��Pj:t�o�W�r?�^�W��R��p��"ZP7����Eh�@		�����,Z�ԭuoY`Y��LF H���$1���ؤ�s�v���Xd���ڝ�u�Ҳ��?��0�k�J4�Rx9��Ӳ�<��ނ��?�ZP_��u8�{'�ݼ�2�9^��$�{�wy贽D���a�6�(-�]�n������Ȋ��&y�[��#��"x.?����ט��C���+�D�?o��5R��y��a�5��.���� �؎jc���V�il�|���4W6�pQ�P��J�j��}aD�ѕ�hhr+,>�Q���e��؅��I�R�f�{��t�q/�%���S-pi�������:bW::�@	�D�9��IU�߻Ɓ|S[�_���
U�5���R���Td�{O�[�R���R��Wds�&�5���A-����ݑ����y�d�!��"��=م7�9��"�����)��	�k%y�
�1z��a)��m
N�=��T���:Ê{2^ ���h���[@0 ٮ�]�9Ǽ��-�T���K4Tyd����{,AN]��27����՟0$ o�A _� �5�Q(����ꂧ�Ir��V��_��drA� k�d��?dK�'�PN���@.Df؟�潻Ɓ�=�'�(-l~��2�H��`#1ۯ�&6����F�7Ad��������ϘV���%����y@*f���.�y�G��Q6R������w�e�̔>�xv�$\���I���;�;�+��1��LZ��f������Ty�*$�L�cj<���wT�b	Z_���竺���C`Ȋ�P~k�M9���i̎O/P��I\#s��5C���;!�ր)���8�(��?5TP�6G
H�1W:5�)0P5e��n{���p<�:��?�37_&iv�6�/�o!*(�^����G��e�e���<v̑PW�]t^*?��.����R�zx���:4
����G/�` ޿�=�)|:������ʣ'd���Lݞ4�%�u��MS,�d�� ���[��*���v{�U�&��4�	��)�X��#�|� [����@2�z�Q���8�⭌�fg����x��f�P1x�{�wпl���j�Ơq����oFF7��x�����q ���*���ņ��	�%��Z�̖_����������כ6�/J�J�����%"���9�b���!��O�-�ǬܚB����Iz����J;�PP�I �fM�>�GZ�X1�_���1<�i�uڈ�� ��-�,� ��.z�-�@'@f�R>�2F�{������9��J�7�zn�l�vEP�*YD.�$���b� ?h����#(֡�o�&������^��|��3ND[������Lʔ/�1d$H��b'�|)r2���{��@5�" S����w�T���v:�	�� ����4��!nڢ�f�ھ�d�ß;Z|>�
��a�0ba�w꿓�XVe�p��$8����5�=��2�"�;S.�ф������F�В*f���?t���"�NG�!e^$ɼ�Y���c�@�T+�s~Ϙ��?.���"?۷�g^�����R�6կ��H�"N���G�P>���.�*/$r1��� �X܂6��O:m+�a��ذ�.6iὝG�S��.�k�i�8$!Q����C�G�W�M(��^e�'|��An�P*bGŦ��p�F�P�(r�S���e���R����~��լ��i���]��Uz
-(?;*=��2r6ֱ�f���:&װ{�3EٓFݧ��/��� &�"�<��la�摙[f<�\t���O���xUa���o|��d�J*'wY?5-�k�����G�9������{_�r�l)/������.���>������������̕��ҁ�Ԇ��Q���>�����mm<��� L�T��hXqKp���5�ja��}���֯F3V�Y�,�kh�i�����ߔ�/Mȯm8#m:����?�=X�k|.d6j4�����Q��+��kcͻM�O�0X����|���C�-���b���l���"'΅��NV̀@�;��s=�jDAMf9.��|J<c#T,� �*����H�^I3�Y�ur�o�Sw�!*���>�.Z���a��'���ľ��cfa0HqdR�`�Z��1���c�#�=C�)���ez���U���#��}�|蝏 ¾�zt�D��O�*M��F\|^���+�F�D-�ٚ��X=��@�p\�u���j�j�eM����}�Oh���2��Hs��;J�2����ʏ?�������&ǥ�n����Ϸ��0=9}o���p�<�d)�_ج�v	c�7z>f~�#����**a���-�LBv�*���lD�9dS��xD�'���k$��r��5��2�� �:K����4�y}z��4_M�Z�}���
�-�������Wo ��� �!�v��_�Ebd����v�;�H����;+Z�����r�n�`�Կ*`>��Ei����h_'�P4�� �	'o��\��GeǍ�*�.[�	�9:C�_s��-A�o�=;Ъ���5$��O�-Ļ��R���~�V�x�Ɓ������6��m��-aS��^��}��{��@Ҁ�㯢fX��ֱ��(�4�o����߷ȩ���y��_ߊŵ�U]��9K�=Wj�����+��7klA���`�O_
F0��W�\:��*�ӅY`��ۣ��f�5?����o�#����IK����=^4�9Z��@�@�r�brZ�1��پ���/�^Y}��̴���f�'�l�'��M�[	f���Y)�^��jw��f]��~d���3��LjE2i��c?Tb>r/�%��cBSM��o�����*D3�}���D%o���[R^Ã�b�3��f�LP��0�;̿�s�X�#��GvS���l�7!��L�qBy�W\$�q�W��Z�YDm>^R��X7�� /�{Յ7�}�b��Ҍ�45f6#/?�ɟn�!3� �S`Z�eZ�t|���R=�����%S�_���y�3�y�j|<����̿(��-��eFAk���
��^�O�q����-��V��[��T|e]��pv��qr���������}�q��11H_���Y{�V�3P�$h����Ó��{�C�<4UWϸ�r~�]�W;xE-�I�GhxN�Z��{]��<�^���>O�
dW�1�0|طa$�N:�_�.6����p�&ˤ���" ��6�,�~���7�Hϼ#�{���\8�����I`�&�BL��T���jB�kz���K�	�I15d���Z�?�y�_����Z���^���V�,nr��W�Us�9�Ԧ�Q�"�7�a�s���=��m����$	8���]­!��)r�W���菛Ϧ=��3.���C��L�;26M� �T�e�v%��yͼPrp"�����޵�;��p�qm�̎<�v�|y����)[�rI��Y�]��Fl��}���0"mcrha�?
�d���/}_,�cX%��C~A9������~�'�[�6ڌ�A�^E�G�c�I�B��A�������Y���M���սk����!�l,��ҁ��G��=NA���Al+3��-��=ɃT��50�<q�EW��>oܗO�=����;��~L�����2Α2�����)��s���@�� z�jmQ~�.�<f�w�}���&g��L�BQ��i�k��qϤ�I�s��ǡ
��1���o������������l�h%l�)g*��5v
/��M-\�Qb��h)�����<��W�KA�ǅ���z�EI�����ڷQ��[G�����vBű�Ap�id�LO�7��O������W8m^@���c_?��锟䳂w1[�ۄ��2h�^yw7���dR�&z_��Z���q�aB֬�'?C������-R�u)��r�Z]�6�'}� lm?aMZ睫�p��MEy�� �v=3�8a�2���M�º�
��K�^�������k�M5��)fw����G��~����9��ϔ�Z�P��f�rUB1��[�W�Ew�`X�SS����}��Zॿk�\��&An$�W��%Ic4�1~~�߀�Gz����>M��!y�������-^���?M��xV��%��U%Ud���6�%#✼V>	pn�i��@�����XXmax��i= ?�Wo��ɰ�<Xg�Sk}�s�"葆�u�8��ʾȘ�+�<�;ں<�}��Q��+\_g�O��b�!�V��#`z:E�E:fμ
��z�&���S��|� ��T�z�%�Hnv -,8Da�l�
O�v.Ԁuo�S����2Y������Ey��N�G<qA	�B	��?o�2���JG9�>b�$OMi�o�+��g;�DK)D�,VF����␼�暅k�_P?�/ID�; ��6S;|8zE}�Q{V�j�j�ك���P��bd��*6z'$Aދ_�F��5�5p�����e�ƦK�����'�\/���&��iB�#��Z,��K�ڑ5�T�|N�-��'������B�a:(���;R� ����<tO�����3 
��ǛK_��6�s�v�z��$G�3�Ze�S�C�8&Vi�Ȣ@�Y����5�������$�}��_]�����7e
\6#堭�Jx8brn��7���<n��pj�D8�̗w� ����e�fv����{f9#ŀ�&�gc�d��of���2C�j,�+^1�P�"X�D�y6�"��{e�S%6oi�Q�1���������>MVT��6�%�5%�F���!�z���k$�h�6J
�,[d}c$�b�VJ-ںia�o�L�.� ���bO�\��j�$l��I��p�ی�f��1��%���J�V`F�FO)P������H���7K�Q�>�w�8
r<��%GɁ��,��#�=�6��WõvT~��^�����s>�����,[�ug�Mw<�t0P�v�|�x�t9�:W���©ㆨ��Am%��p��O�r��n7�j�懼A�Ͳ�;:�&:^T�#��L�d8x�>�"��$�Ί!��H�N�Oo5�0�꓂�X4��0����6�j@r�!�Ȼ?iD�.�~	ҪLX���uٽ��ű�-�Ⲕnl�dÊu؁G�Ts����=i8�b�἞�n�y�D�N1~_���ӭBj+~�b\M�8 �4'�m��ޏ�i�z�a�a��@Ĺ�K0Xo=p���GW�t�y�B[�Y��Co�H�e��5�@(j_E�R��QO���)��ux��pކ�햃��
�wN��/J���N�����9�%�����l	<�G��Z�L�\�I�76;�U�� xsȃ���wɎ�-�]9)�ڎ>@�H�]�(~��}^��X.�_��P��<��˗*�,�B���L`��={�m4iο����3р.��N�@�:�K�#��ݣ�`ͪC���m����D��E}�ܝi*��z�B�Q���3�@��/�*8��*�H�13��m�����9��)�����2�Sx.�l�?�Qhƌ�f;�����V-��l�?�n(�� ��mz��,�=��Q���|-�j��}�����(�	�`{S������[�+ ���B5����� Ȋ4]HͶ0M�z�P!h�_Mp �����j�My}��(O%�p.p�DSK��L��b`n�\}��� �pL^�9L�'�~|�j�ʌc����J!4U�ZK�`����A܊^�v����Q-���C Y巧\��*+=��B������U��`6#��CF]�&�O[$��s�i��T0�*�{E6���k���*IMSF0�)�����J��a�$��SÇGUۏ�������wP��Xde�ޡ�s+0 R���t�	���m���t�O�}y�
�Aavi���V�	3�(>��}�CYtp�R"nϵ2�l&4�q`�J���V FwV�ɋ�̃���|}����h�H�^�pŞ����3 |lW(�J�(�vϟB��	�뵏g�18n�M�ly$)��(�ys�|��k��}����q���Q�W�_�� �Yb˱hY�D����:w� �%϶w��;J��G;�k��T5H�9�U0�spiW���4�]2���疦���r�x�|��0�,�j�E�}T0�Q�x@��\�7jQ�)o������ۄ�(2 j"�&��}�lZ�|?u6F�(0B��/��3�O��<Ɍ�:���a�v�v�b��4\�mpK�^��	���Yo�0���B�r��f��Z��+��;����Di�FeP����2j�^S�:ޡ&�Bsػ�foXmȯ�֖�.�=�x���K�"�#�x�O��&�4|�!q��0|���5�
w��1��g�6�o2E��y7J&q� P�G����/H� -n���F�.k=��+�§�t��ub�%5���v8��L����S�jTf�}�d�}�P�Wu��'#J�9�W�֕)��s��{�݆F�-�� k
�Jř���aN�@8H�^۷CVO5UK�`�o<
U×�Y������C���l��˳>�L�O-���D�����Q�.�ںC��G��q�jֵ�m ���;Eҙ�0F8M���{���7Zu�?o�'z���Q�� �Rm����]0֊�E� Eq}j������W`�Ɣ �7t%h��VC�����h�g�VAJuD�~8޿fq"�ν(i�� G��_��q�A�>��� �vv�J�5&(<���z�fll�:�}Kl�Q���RJ�VF8I��H���@�w��t��ov��\���[�Ӧ��#LH���,L~��T	Z0!y�m8/����s!&��m��>x�y�mn����S Qr|��,dܼ�=<!�7�Ye��ܞ�%̡�Ocm�*H�^�LZ�:��#5�M`g�{��t$F'���qL9�.���/mla��f5�ݱ^�Z��K���K2}Z]�YI������ܼ��jt�ou��8��+����q1�C���huW��mA���8VV��wF���X����M����j����#����1��3;O���x�/�"_p�А�L�&����'�dب���c݂�Q��t�Pmw��ݳ�K}��Ĳ�c6��NV;UGe�M\�{�d+�P�n_�[����0���^ꙑx�>i���T[5�">���r�A��m!k��α�� ����kFx��/��[7.�
?̆'Qf�@߲mE�Rupf9Ås�b��@:YHE��>��x�&|�V�o����9�a4K�htw�����
B	�3��;���=��%��1��/�'�{���o���D��K��>�ޟ�J��Ύ	�I�r!d�I�y"� �/�[���xݲ�r]���b����Mw+��p����]<0��}��Ǚw�@&��4�.�iψ���/��!yD�.���:(�c|��F���r7H�i`c�X ��@�����Ε�S�C8p[��qy�4�?���j84���<b�G�����랦.�b���K���!�`�By<k*���0ݓ�awěF��^an�;ۊ����{(���@��h�߱�?�jk{7*z�u����XI
�2�~��{�ˁ\�S'B:j&ΒlM���s�ӫ������٣>����5>YBY{<�0� �6�x�b锎J d�N�@c��3  �Ͳˉhu7?s��-P��v&��EsJF��$�Z�H���腰j����b�6K�(�F�#s��ǲ�Nzit��~q�&L��+�ˋ�KL+���H��P��<qe.��Sl���$��hN�W�!��
�ר�18W�{��i#K�=	�7Ԇ+�g/�h >�t�0��={���R����AC{<�L?�!��;�kE
�H��+en���kS
�Bi����B�#icH���WR��4D�S�#���DX�Z�L(���D��#<��ÿ��N�(H�"��� �5F4�D9�>�l� 	�4!-�����x��,s�d�n� ���ܲ�n"$��d�#�|���荭c��yujh$���^a���q�ĬX�~��/�������$�*���X(�h\z2է��'M+@̓��a�ܤ���g����]KD��ϴ�P�jy	��LD���;aq�Y��������ϙ����?�ġ�MUZe�D
�
�s��D���T:�d^��O��r���2����L��4S��O�����}u��NC��Ⱥ�����voP�#��н�;�B<�M�x���B�
V��R�W�)�[���՞ŀ�==�Ј�&4 h�/����W�����'�[{bMW]W�������6f�<�q�s� �k�0W�)��{�����P�rSc��Nq��{r_�^��Nl)�n`��v�ȿ�␮VC�LYb����&+�,��2���A�&*�����-, �ƣ�Leof=&�!�#�i�y�bn����8������|��~e!����^R�;9JX�&i	��U}�[����<�'\`6��4_�3a�wz��� ���H�6��S��^�VܯU"ն�`�:��䩉��i�bYb	�Z��<�B�����Sq��*1'��7�c\Y�|W��S���G�����˼��s�����s�+�L815U`~��-�H�A�0ʁ�%����(����b���Ŀ%(�$�]�O#yG��av6B�°��W�Sg��!k��Y�75g����+^���_�}��Y�)p�M#�l2��D������[ke��JZC^���C�e��v�����.{��J�sI�4:=�� ��2��`O��F�{Q�m�KjW@x����cS{�h����03>�&%�3��Eͺ5�^���}��Z�ZϘ�)5O����=�:�ަ���|��4����\��+�1"����o?%�.��]�wb�VP�C�z�0.�ڢ)���͂��������WX���a�3aAd��M�zԉ��������Y�P��S�<wr9&��:����A(@��lF�;E���2���8q�P���4ʄ��c[t�V2�C�� ����RK~�mJ��F����������5�a19�q���Ҕ��yv�JP+y`�c�hY���њV�}q�ߌE�������tjq� .�V15���N��鸳��%;ӆȇ����8�<�&6p7�^�f���R�ƫ��D�������8��-�:�z��!�^D�A�K��P�##�7F���p�p5������82v��`SyA�t���I^�gsa���#RٔB�`ןI)��*�����f�;`T�|�x.}3�1���wmn�j�§�wv�ӵ����wB|��B�������ԐF��j�f��I�Ўl_`��x~���0?����u�Y �BJ�ْ�x;e\�Q��?1�DԳDЊ�����G��~��~/G��18g��R���%g/�q%O�L�tN ��<3��y,��S�Kis���?	D����%��d�'��I�CT�ǡ�@W�ܰ�\��C\����;���ss@�d��.>z���f�����`te��d7cݛ�̚�A/��=R��3%߃��'e�p���e�@��2#3�4��x	��~��v�i`%Y�	b�n��9�b��.��UW��1��L�ː�Ǧ�&�ga�H_�Ș�tR��@�y�@׷�Y蠮��K�0���.Xa̝m�������c�n�̀��L�	W3һ4D���Ϧ{������?���*j����w��`�5���R������❳Ō�s�:�J,�֯���ëӡ�<h�:w�7]R�^7x8���:�2���֔��դ�Ǌ$y�A����@<v�����(����� >
�b�P�n�~����� "s	���IIHV��K֚�:�|����B�� �J6��>�'��k`���.������!�P21,�$����-k�r�u�8����D_}���1��.݄��	�T�T���,Gk�-��q��q�s��S~Ҏ�+���0�;���7���s�=�.k��\�.��.�kOY�y�y���HVN�qO��v �]����@�i_نi�vQ�bV���j����'Q%��x��mkq������"?86����!
G���{�F�B���_�	d}0`n�W�CFY+t�/�qE|:G6M�{���h�j�â�ݰ6�!�ٺ�NG�����3b�Y�������r�i�c~�&x�+&�:���@��ͮ����}���k:�`�W_�~Bߘ�O���Rz���Q�q.`�wU^'=5�4z���rlA;�Bl�i�c�����'V�|'�b^�H�nI�m��Ԡu�-��8K7Eg�'�,g�K�䴭/�js$b��|�����D*]N7�P~"�X}�eh�?έ���J[� �h�æ���c���)��T�e����P��A�Y1�� �<ů����o\^%�Ք���G�6�u�G������G�|�@�:F�!�)��/�Zi��7�G��K��g�`��@^e��~�9v���f*��xYn����)���
�ڬ϶3M���g�d�]�PL�&�)�t��8 3�?pR;y��c?�utYя��]:8w|���&B^e^���rq���zU����
/����	����\N��NF�G�p��3��'�I9�8���]�1S����l�v/�c�!8�q���� ��8&�#��d�IL���\�^ۤ�����mn?^w�D��]�6F�x�{��Hk��O�7ţ�-�s[������'bn�(@]��(�P���p����x,�	��:4g����7�_t��mÚ��i_|�	A񁕚%���i	�>�g~��e^'$��^��1,��>'W2,��)pĕd,��>F%�k��2�8�K�o-'	�p����0l�/��̔o�woۀc�{����H�+��ǽ�{h�?�\r.E'���2`��u$]w)���H���8%��4���A3X���_2�(���A9?x�8+��d�%S�2N{���۩�0�� ��߶~r>K>�۷柪#k�UF>�ܭ�}8�A�s��r�<�G��Y�j��B��s���,#���~�>���^̷7%����;�g,nS�\�(�ڢqjƓ�m��k��?���AC����fOR��th���T--S�P�/��/�M�Jˁ�䊦�/#�4*�>w&b�	��~گ�Ef+�t�q{�>�'ؑ�4�?��E|�[�	�L�� /����R��Ƿ�ĕ��3es�\�x����<���`S�`�s0�M*:�9�0�F�*�͠[�]D�&��^	Y�8_��So�=]ˁ��k��l���@�{}P��3�V���9A�ؕ|�z��H';V�3t Y��5���7���ʶ��O��z��dmR�kc���\���� ��+�r�V)q���\ ��8M،�:Ist��S`Ѿ��ѕ�?�kI���;54d��w)3v���r�=#���S����W��2a�턓�B.���(� -�����*}���|w�5��kMe��/�'�?���H����F��^&�'?�ne�X�}��)�ԼIW���X��a  !l"6w����� Q;��d��^8m=�g�h�24!��u�'�j����Ӡ�� ��:�u=�w^=;b=u��>�Ӿ���^����v ��p���Pp�����S���W�xpC�n��΢\, MB�Xx�&�å�F0y�(��1#����l�yH=�Y6��?`:-�T�.��@v�l�Nɟ!pk ��l`�2vC	�����{�|h�3a�oF7Ly�m��D ŹAC�Ί�U�T	�n*����/���e3�{�H[�\�>vN�(K!'�s���!v{���H���k�K"A�@���f��_Ocƒb����&��ۨ\=��e_@X'����I��'a0J��,]�He�J�S��<���ϫ��;H�"��^�Ү�r��3Hi�%���(�\���٭QN~���oWu�r�W^v�� 3"U�2��w�P?�9ד�o��[�r�v������y�^V�f${�Z���MG�Es]~����B!7i����Õ�]�!�f�
��F� o�~�6����H�k��F��T��w�$I��d�$�n����ғ,����eM�.�Q�<���G�,�1�m0�cE	F���E���a�>��P�*e�S�|~�>]d�\����p�QJ b�
���-�����O.K��	֧��Ѓ���O�/�l��Z�l��C�h1?���K�z�\�nS��'�KUM}�K���e��t�$�C���+�?�J
�70��\aѓEK�5���Ֆ��R��g|��� ��/�9A�0�v�$��jlV�E!iCz]D_�UG�AxV��m�	̅�;�M')�k��{c�;r�mQ����c����������̎���{�����G��9.����%�Y�qH�Fo�U`�g��-X�K����JE*�������f��4�P��j꫑q�IgG����]^Tf;���smo�Z(�=%g��Db�1,Ma��so��
��ݴr�:��������7�{$<-+��t��� �ק��K�"l�0 %1���"'�u]#9!+�ؒ?�G�Jh���j?x`���G*�*�AU,�2��AF�_�At�Z�c��U����Y~�Oq�J����2:n����W�ÿ��?��� ���:	�_E���$��,j5�fcK�'&m���L)�O��J�H�:�Oq���/�l���>�0WǄ��	]j���0:���y8���ԯ�!ja����q�R���͙նho_�:����z��7�~�&�4��Hg�����I��h��p�t��� 2M�B�VII{,=X&�R��i/'v�0����P
�^{��k �iݼr�rEf�i�V`ާ���m
����kp��y�$���Y@�@)i�'K:�G"8jZ��f�pY����>Y�*��ď��N�.�U� �X�N)8qP��66�O�AK���u��u��*!:�ǰx󁛸���C��>C���p�I��yG=��iM�\7I��U�8�9m׎I�^��O�	G&�ԥ+D奎?%��ŔkrULW>P���},0�DLq@��g��`5��褲 ��luÖk�sW����P��F�p�$�.�W/R$\\��6c���p��f	��0m@<-���v�c��:����/�D��9m��3��wi�3 ��%y�h3�����ù��[}���7N�c~N�1P�v��K�殇6׆2��I�q�"����R's��^J\��9�����y�R�qD��j�҃������N
���N�����8)5��J��Ǣ�f�@��$�Ũd��%��h�ٿV�
�zs�M���:l���3�d��J�?���sI���O�o�z WI^@���B<U��e���'+��'��{\rFU|��=���̖yn
ӕ6.?Q��1]�b�p�1��r��*"/&M���f��+E� ���p�X��0�*1-ܛ���_|p`�T9.�Si�K��km���)�����Ԍ�20[���+A��h��V] �bi�;���+�)������ZE8'���4ػ`PPȆι�r����#7h�3�*�!������;W��ߖ|x��sQ[	��6�1G`-���;���7A8�$�c�ǘ�YF3?ݞ@�X�;��O8G#�"=arw��{�^��ܐ��e�O%��K����3����9wauh���$r��,���V\�gE�С�as|�T����!;�+�gX������v���SP*413H�z0qyB��t����m�C/��Qx~=Ma"vJ1k��	E�D�bu`�~�?����	����a�x�ݿ�S̢Kw�@��0���e׽��U�<"Mm5�)O�|O(�dyN�}A�fm-�8�8�ĝ?Z3��}~sѴn8�K�|k�T9!�/��9$��-h�����{�o��'�!�I�F� }t\	�m�"�B��8k%S��*5����ܵ^i��8ԷoT�����O'@��ńG��PgT�ޫ^�
��5�2J9��%��Ʌ{�[ժh�?hę����{yQ��lZ+��vNp��u��*=eI��	g�����i��ї� �Kn�ӡ���Z�)�~��#��dn��H���S}��)��]&s���e�H�wn��2鑗V��2�$���kU��6���=Q��0ڂj�_��a9��﫳#7��;{O�������i\�gL��g}�L�J��Y�Z[��l9��{����C߷@7�����~>�TA
��M=A����ef�+����<� N��/�$��{*�fR-�����r�`��W���i�ok�ۚ����[�`�s/?<�]�F*�Zj��;9x��[����B�u�����-_=ܸpMYB���^cP68�@+�[D�`�rdR]}�iu�����uxd%wB׽�hf�M�`�sd;��џ����B��<\�@�N��om>����ݝ�S����P)�B�[S��Xg�b*��׎ȹ]EZ�2#�>�^�$�@hhG�+t�c������,����A�� �W��h��'Wg��%�	�������Ǣ�Yӛ�mQ6o �u�i��&)���T��G"	�̭e��'�(��^cI������FLE��P����r�u�KAR�U��bl��s��J�5S���r�@~�h/j��l�	]$|��1{61[f�Օ���X�h�;��ª�xj�6D�� �	�����`J���K�f���^=�@�FX���X&�Y�2�Ns���ۂ�Ɒ=�N��v��:]d�,��<b��u�B�r�#{
=i �X�NX�V���������}�Zq4N��[(ݵ�hhR���O
�����g+S��F-����Ƽ3�JX�W�Q^(�+�k���	H�ɯ�3��3��u����e�F@��{��N���@�?�x�~��%3��ks8� 'f�+�FkX�]qr�"�',��ﱹ��XK@b�v�(�È�̆G�X�L��qsǝW�v�WX�<���nX��� А<�*sz��#�#Mhw1r�����7}�F������V��%߬�|���I0\A��Ѡ��A2�̪�����dj.�$������^�᝺C0�.0n)F�����HC ������|��51���k��<�"#=�C��9���lC,��`����m�S#v��d�,�@��퇺�i�h��1�������$�@{���e�T��1�֌Ϧ�K#py���zm�?�7���߰�i"-j(�3�6x���������3���7LFn���Q����G��ƒimP\'����J��[zɿ�!8�c|�A>y��❰�̷\��gnU�hi_h�
��(*33����V��D�r	��,��k��n�� (힔
���s����P�݃��o������Қ>q�+I�OHwu�����B�Toz6c)��`:�?0�g	`g�ZO)%���+0}���ҸH�g��R0��H\ݺ!1���}	^�=��ۭ��K��ⶲ��_.i��\��&��	1c��c6�O`�_���젛ll���Xm�)���&~�s7IZ�Y8�3��h�I���o�l��%���n���|0�a.Dp���#P�Y{�C� =��� Knԣ2�"�+n�0
�щIh�F�Xh���8/(Q����9a���wvg�P<p�!Ċ۰N#��\~N���]�	Z}?Eؔl��;�LK0��Ѽ�1I��~�'p���݅X3�� �b�o��M]M��Y�& ������kO��?��7���jf��3��+���C��܀�p�[����Ň8�,��:'q�P���Z�,J)�2B=:��	�H-�D7)Sw#������.t��]��Ζ�|Hr�g���U8fɨ�e����S�3w��׏�RG7��Q�]:e�|�J	��Le��1���Dbrt��/&�s��ai��XM/j�2�����~r�ʇ����+2���ք65h9*/��6�~��� #L�혻�JY��컁#Ĵ����K����M��������I �5;_lm\���ay��!fR�� ��T<7*�:�J��p2��'��6���7�MF��}�r��Z��3���3J�Tg��_.=��nGI\_Ś6��f�{����Sp̒�EH~[�t&@I�oED��qჺ�C�_�!V��2I�u��|i4��I�,&��#�J*Bl��?� ����Xp��-�ʨh�V�pQ6�.�O�����,'h��D*�@�{�50��LϾ"w��?':�FB��S���>c�)=��L��
Vā8=�Ζ
�X���u<X����@���7�IPӚ��_'X�ܹRY7��*FG�q�6G��V[D��|4���&}��f"l��w�f��wӅ�I�p�%��������YL�>��Do���#�#L�mm~��SԨ,�1�&�;Ha�r�]��j�f���� pk>�0BqK��oF$P�[5[��"��pR��/��%�!�(-��5}.�~�#�Ǩ-u�J�k�˪c��ӵ��[!z���27�}ʟ�t�(�X��9�l��+X��!�=�oU���q�����`j�����O���EbΔA�۞<!�����S�R�W7�����cd��Dih<#��L�#������x"���D�gW�|FQ,��q�]��ƀ���(�]�SJ��,�PE�������gs��%�w���M��e�+�.r���[�@d�
�O0�z�E��u�0-�d�t���~���>��5�x=?�6@�:��=x�z_�zӾ^�2.!^�1Єb���q��PvN�0ޚ��=q%n�a�E+�<�,��60��+w�!�='�{q����|b�1�%0�'����acJQv9��?�؅�+�@���_�������r��=�p��`C�N�Ż�4t�ԅ��%+`@@��W#.�{�Lb�a�#�s���
�����~�IP�$\ �6�C銯�!�\���Y:ɀ�RX�"j20������y�R,*{����j�\8n"��m��v\����*�Ag�?�v�q4�|����]s�B����d���$V�8���6̕�����G̳%���䍻R8)\p
�������sj����)����n�a׳E�M��������z&!�@��|�����e�����;z�e�;����U;F�[���d�(A5���)�-J�ڥd|Ä��ݾN&;��4�Yx��-_��!\���[c` 6�V��� 4ߕ~��AK`��dU�_�=dXw��}$u܊37�1�g�>M7x�O��D�3u]'�����u�*DzM��M۷z:�G;_��z�B������;̎�=+�D��7 -Fø��x�q���/9=�l��Ô�3�m��Y�-��Zkr�J� �A1��T���,�����`����)�U������sN>O'��}��2IxRy�l��8Y��ۍ�=k��!���8w�֧����p��g9RÙ	.����-�m�^�j�m65a�����A�)��]m{q������G���t5�0��XE�]hS��o<<��ӉdAc��/�z^H	=��Y�Sܞ�cC�W��j9�Ew����:o��{��O���t�7
_�Z�x~��,���D�_,	�^��]�)�Em<d"�$Sz;�;��I�j��*�_t$�HD�+�m���K�B��d�(������1�~$9�z ��,�ԣ�z�o��x���-��.���v�gI��X�C�0���C7��W��qZ��y5�@�~9�@Jk��U?�r���|�L���e(p�wU��?���L�G`Qla'�\��dkz߆|�R=�6x�g��\��G5�4�m��?-i��xG@���<�8�a';�5k%���]Q�Ͼ������|�zt �:�T;\�����\���Q�@z=�a���Z]p��^z�.��pY];�x�ZbV�f �G�_ߐ�(F	���E[�|ޯ��{�U6�Q��0f1�*EuUM��� 1�����?R�H�2��SN�n.h����? `��3|��^�oR�ϱ���w�Q� ��&��d.)Yģ�49��|e�Kg$O�m��Xdk3uȪ#sU�]�8�cv����*� LJ�a�oQ�\����js���:_��q��o� 1���o���L�6}�h�щ�=��?"B~n��d��>*�30V
��!VE��<`@�񔤴�M�q����^`��i	J�=@1�ס��I��'���T�*�W����!,�� �^��̨���d!�v��#T��~�W��R�+�0g�0�X���񲂒)v�^��vw'X
�٪�؛-�Y��A_�v_E�E��0�*�" o/��H�$$b�
[4��`��lF��jy��x�_��8JC�?"�.�g`�?����a�[Z����;aWuh��EqN1zvR�9^���P�������nW���ɹV����6��	uu%����m^͢��{'< �ѩ�l,�l���Mc�R�*��U��B�lЬ)%uw�ꨢ�FQ[e��+�Q�^S���С��x4|�@�nX�R_������~���]p���&��a�8��Q��HZ���Ge��%X`��oŞf��<W�?�\��!�v��@�hU���U�����יR҇�P�x��<�����ޙ�L�t%����������M8`�a��� ��`��`�xTǧ6lDp�H�N�!"�.~�Uy�_�UW�ú2���RQ��o�,u>{����PT]��V�]�x}�-�
���1ɬl�B�������9hgM�Ø���-��Y{��`о}	�/��uNTxd��};�I,J�tuW��B*7!?اF[�M�(\��h��Az�@ZAR�	�kf�4�����_�	���[�0f�������T	1	�a���h@݊!%�.~���2��<��ݡr��b����<���x�U��٭�]��V9T���}Y��Ԭ�DX�o��K貴�!2���-��ި�e��F�t�X[�ԇhֱd>!	���������L��3��aL��^��5]�n�"AO��=���?���Xbok]��1>ܤ!b-��V0�g��v��o[Ӄ�p��^0Y�o������O�fI0�+Z+۳�`.W�x�:S��"C o|�k�f�n�ܾxͤ�'�.�wTmjpWY@^v�ōǰ��j�Sv֋�hK��Y8w�Flְ(��::��I[5_��0��Wd�zg�:�fJ$�fB�਑z(�;	^�t����&��H�l�bO���.y%wH]���)���?boT����s���zdէẼ}��C$�/�Ql�F��z��
���w(;k��.�c��(��=�_�Y%��1�W��t8'��k���kFUc�L~���
��%��j4���_�
�n��P~��M�6���^s��a�7Rv�T���c���)�j�)
/̸WfP�����Dt@�Rh��9�;�3vX�`����(��*D�,�so������G%�n���;d�6�.0k� ~��'�\�m���}i4A���LHJ�0;���!��x� �ԑ�H����wY<���?�(~����X����vu���T� �?��&���i��e�=@�Ӹ+ȵT�ʧ�M�͔`q�{�y�LˈS-�1Y����L�J�#NX=z�۷jmm���o������*����Wv*�O����{W�+P$Ã��*FꠧD������ �(VMk�P���(h@ܻ�s�Ƣ콟�(��d#E1��N�f�/�̲�F�8���a��R���E�#Ｈ��ڿ@�kD�(9�Q��#_2prϾa[^�� �Ө�� Ґ��"����$վ5eQJ���Ó<�V:�o!��L�V�l!)n+xI�P��q�e/|?(�%�}��8�������l�pI��F�y�j-U	���<I����H�F��ۉ �$�0�6�}u�@�v%�Z�2AY�B��|f�hC5^Ca0L8!>�����(�8�?닕|d��e���Ц��u.���*��1����&�m��<�,w�BӸ���9��
��S��iҟn�Q�����C< /��T��� HND]���3��ee��f����] A���~Y�{U�`����ޗ.�_���b7��t>/QS.���m��Jq.m��r
��552$l;�'3[̸N��.;��l��鑸�b��g��0�ު��7��i�oj���
������4o^WOt-K��� �iI�t�uRGR~{�!��e���ɬH5;,�j>yq	6�Oj����˨;��n$�`���I�9k�%�u�G�����/R����:�������=>�
��9��x������L74MS{+�,/Y��:�ߦ��P��V�dӤkJ�w�t� 	E���;>{ �����,�μ��%&>6'n�s��G|�)�&?�-����Qb�^S��/��_\��]��*����/.;�|(����nʽ��<p�4�'8��╃q:����CC����s��a�����se�2z��~YJ�2P�G	erp,|�,�����zκ�Џf�K��W%7EL K��Y����WfV���	Ve���K�s��Fㆠ�1?�Ӣj�'�m�]�	vb���r�}�F�FԚ�[���R'�Q`XcH##?��0u��U`3�idJ�성��f����P�CN��m��T.��*g��<l��	x`<��s�"���~V��"5<�
)і�"N��_Ӊ�x���	�ŒO7+�=��j�7�}�QuHb0{�N�T�􀣙�6�0䟐@��p���"|�B( ��)k�P�s�|mA��p���Jlu��UaC����fG���������w�V�(r��[��l!�#��"CNOVq�ȶ'�(�9����K^��:�[mdY���<�(�(�1*ַŵ��mu���R#�7Xz� �?��f��߃��l�r��hc���r���Rݗc�Ƈ*BUX�QC, �g���@���M���%/ K�a\o��ƪ�p�	�:~�=�
@���]wc@�~$��c���%|�:dKPD}r���Fm�xe��H��g��Kjw���_�1I�|��Ob١���aJ*ȃ�b�FB/&��L���d�_�_FEN�g�Xq�Ѧf�q�}[m�fO�YS�R������%;��9�6���^�:Ș�K�K��Q�$�OU��Z] ����Z�=�$t�1�Iu�z�:�w�_��e�M^'�ѽ3�Z<'t�ȍ���y�OU\�V?S�<���o��$X'��$����fb�m+ϟ�׭�B�?R��H=J�Ыn�����oqi���>�6x/Ep��fp���YO��Y˞�E��w�b#yT?���Wb5N7�L�&Z-<�BK���/R� 0���=O�P�h�>���l�1~�� �P�?���mTI2=��FI0��q�:�Zz���� �M�o@y2&����E4ľ�x��^3v���M��������������Gϴ8T�M����ͧ*��Zn��j0w�Uufc8�b������N� ����A^���Y���@�A����ӏ�G�Ꙧ�9�������mKOO���n���w��������א��9���W��w�f�P���e���O�zn�y�58m���^�q��\I @{fQN0(F'إ� 	ţL��C�?�N����QD�"�uÅ�;�EՎ֍.�jI: #�܌�nk�|y���Bo�Ο��xő	�4埉~�kۗ7l?�⩨cC'T�[�J!�Ui��n��0�S�p,`V;���_�b�F�!F-�\+m��g���r}.���������n�+�,��ֶ����c��x?�28��E�Ҥ������r�c�皇)��y�$��XP~�l5-IN~p��?a�S�㓘��D��vj�8�<j/+������g����m	�N�g����I�ؤ��������E�Ѱ�73���4�d�Uj!���ݫ=bF�=���M�N!��g݈��Ȇ	U]��SS�P��f�vF��=�g$Ga��j�$�f��2Wi)�e�o�D�r��Ȇ��%�QM ����VgTY���H���m�;�EȦ=�%��Q5L:�����K��fԮ��bd�.U������b���1?�؍�7a�8�F��s� ��>�I�H�*�N�=���َ�qA��u�4\��qE֐/q�L���7h�c'c�߳ӂx(�~�'|�H2[�P>���m���Y.�E>+�Q���e{�n�'D�ǣ"fE���$4,�%JMd	���t6��Ql��(�q�ʷ�HG�e�By�����QWa�Y�����ńY�����r�����3'Yf�Eo��6EJ���|���Q1?e�V���f�}����@e�5�]h�FCc�)Pb�RU�겑����l�Z��V3�F�T���֔ʥҩ�K��`�ߓ-�������=����5X��Ƈc1A��*��aɪ�L�2˅�
I_�b܂կ�q�-�inlkZ��*&sA�Q���f��M�0����p(�����\+��<kXv�eB�r���6���E2EX|�6��o"g���Z�Ʃ�?���'������c�H��rXv�4!8��/�r��Sm�e�]"�-v�Kp�����o��2V����uPf�gs\�E2{��d6|��0�ۼI�u��␟a��"��k\o�;=�,��r�P�1ٷ���p�6y�Z"�ԕ1?���%�d�,����'����1�a�'Pv>�SO8h�3�!�S�=��+�J���B�!��@�C�;MA�=�H�-��k�/�v�ü��s�<�)�:ə��{�M��=��I�~��Ї��_j�J���!�8�M�j�v-��4`D>���_����ss�ET�Y�J�K�W������;�>t!��U�O?���uq;��T�?c����o�k�\���. rv{�J!��[�e���[��s�F�y��٥Zs.4�A?�+Ϻɴ
&�VZXb�f�>��! ��q�	&���V	3�(,�n]"`Զ0�v���b@,�-��9Q	��^�@bz��Ϋ��8�6�|ݏ��?�VJ�1%T�ہ������28����)�Q�ZQHE�~�{�\�9��xy����{C��������}� sRۄ<�û����DiW���Zi�ܝ��؉U�����r�*� b_�Ѧe�-��o�M#c��QV�>V�,%e�=�u�aku���L4�.%Y��8	ZvYx�q0��hK�dV-h�?8$��w�·����P�3�|����JOyy�SNn�w��f��i���zC�P���e
�L�.K�`��O�o.��y�j�c�}���0�Yu��*��)�W�|�
F��VX���$�Y�[2�J������Yc6�o�={�$Ƕ�$t�~'	�b�\Q`bÕ��8�y��w�Y�{d��t���c���{��V��mS̘}ۣ6���O�5���@�b��0�V�+�\�:X���UW�jR~��̡�x`{����a>����6�_���q�4��"Q��,\v�z�@%v�'(
a�x�-��p�]����v�>��G�b�f���<��+YcnB��
,5'Y�:�w	�c@�xS[C~MM6�h펺I/x�WЇ`���o��_�����1C>m`�Y���N�l��I�sr��J�F�����EN֝3~/0ݗ��/@�N���ME���2��X!�D��A$8��2\v���͎B�����}A�j���9�x]'��g4�G�}o\��OQbH��_�GF/1!���{u��
�K�TC��@t��ۂ���E/��"�M�Fl�D�8�N4�FR���g�cC���R�Ĉ3}& �\��)K�1�7�o)/�My�����"�Jm��9��0�A(��cQc�7���}lK�`���z�a#��=d�!�a��M�a����T*/p�%+������m�Y�@�_����q�K��Z !���/�Pf�1�m-����F28��Թ�B�(�� e��6��[��(��B<�!n5�rp�~$��;/) ;�͡�L��s��es���S�c�P�q-#Nz� �tؓ��g�*�i֍c�;����f����^o�SL�0�qd����m��^�/�"4�@T;��I����X�zN�w,�R<	�:xʅlƦ>3�r��$�mv2��e����~@$Uf0�O
r[�kU2�v�E�����1Uu�1e_��Ջ��E^)�����}���a8����+�����'�ɳ�vUL՝�F���3�}�*ی�!�G�[P<P�L�N�A��.�BX���@�< b;d����A�ܱ�}�n��,��߅?���}6L��h�߱ue�Op���l���b���s�g�5���I��h�<������zb�O�<yQ�Kisy���ŕ6w���7��1�aǗ�c��� 5Y3R=��ݪ����iz&-ԇ��#�v�y-Գ��U�D�E�?<Z�����􉠃]�F;g͘p��xbpظ��Z�A�����gh�ݦ���.Ƹ�YT��z���ɁG?1��h�W�U6�Â~Mz޲�]��M�B���\_3�~���<�3�4��6x�/��?k�Pu�G�˹2a}��#�/P�f��g�/�B��R�"W\I�:u`:˒��k�7��ql�K����l0JIDiR��1���G_!���~UjS����*3.uZ}�f��4I|y����ٜA��,b���Y��6�"��#'���$���LS�*$��`�=[�0��w*�@:��T�$�n��yT��\A�	;���eذ~�X�)������-�!����ݲD�-��qpF~�ܔ&��]��J�/�<��0*#���\=ao��rǻ��X�u�f�����7�L�����9R˽��(��r�5:穣� h=S6/X�7�Fv�|¬̷ �����%�]�=Y-t����I{��)�`�_�];	�"�4))�ȎP"�����uI��=b�	��`'�w�EH�|��������P+Ky��ʲˡx�Z�z��֭��ACPe�-�(�����L�/���J��+�+X��&;1$3��4���1�d1��ż��=I(��.R�7ŏg �>"{�}�V��+:�m�\L��rJoa)X�f2�9����9�? �yg"�pc��^�(�T��8�K^�Lsl���=��|B`�dSS�.ߝ��������ؕ��Z�/����Gp�"쟜�p��C$-kl�h�F\|��'��Х{�1
+���CŖ�Q2Є8ך?M��
v4�V�b���%�m�lY�n������0,�I7%�5B�2J��&�c��?h�?����Sgt��`�������e��F9Os̎�����捼��E��� 1�A����a�m\�����EHq,���L�}�����<S\��!���*��o���ZZ�+[�s�1a��n�|5���a��%=j�΀C3�8�Ё�����>E/�N��6fO<k�z@���Q�-�T�m�/M{����Ly�"�j��T��o�^t��/	���R�p��/�r�n��r����6Hk��3�j[��x��Z��1ؼ1]�T
��6*�cf���C|�9��zk'�2{h$�=r��k��0��.i���������'�zz0?�aZ�4��_c~��Hw�WmBǱ�J�̣�F�D9�'�\l��ń�e̤ԣQ.��e�oJK¿��FV�����NU�"�R����^�癗�$Z�-�'��Ij:�I�ʳ�}Lʙ�4y��D���W��x_���蠝s�?�q�c%�AMN��R�#%j�)��|h�?��v�ku�;� T��r� b���+Hj{�_�\jOo����u�"����;kѬ�<ٞv���������݈d�j��9hz����U�5E�}y�>�x�>�]��>3�uu"�ou	���wK]F���A�ݯ��������$��r��} a2��ruC�OTyֺ8w�&<��9D��4q��aA����b�j�X��&���"��,��׈��n��� P���<����[��ޗ7�or��,|,@��'dEŌ����5G��� ����j)zr�:R(}�[3��42�v{�hyX���V��{j������A��]�Q�j܃d�!�}�o��]� E[�LW� �*��Hݧ �P�H/m�@�M)2�z:l�:ha����4�e��\�1lJ�󵢗�M�z�c%�u�����e_�y ����|��f�:n����_z�]>�6��,�g�B@Xa(vq,׫��i4�u-����H�1o�D�d���O<߱�27�)`���R���Z�;?��ءt�G�v�BFQ�������թ��j-�G��:7���?��o}�SL��@q�(;<��J�p`ό�b<v�t�Drg�y��&��M��� i��ؿ.�l��7�R��#�����/�*'��p1���U�͜o
�Q��eeyb��0�M����>}�jU��[��a�Y%�a�̀y]�E�B[����7��Y�=��,:��1��̧z&�J��l�m���Bq���A$���EWޚ�nU=͎���3���>�^ 6�i�)�c��d��
��pK��P��ZuD��3ǂ�y2�v�fl�x�v]�[}Z�ϊ_q Ҡ�S�Hi��'L�6��я�*JRC�%q �Ǎ��$C���Iep�ph�f�p2�+T���*�����&��G]9fKq�,e�)���0.Bɛ��}��q�\ؤ���\���7ټ�'�B�)-�E�!?�LA�H����+F^E�̙���׮� ��Y��U.�D���_��{Y��[��i�T?U�{"��USG3Znp�fDY1C#������>w%ը��}X������/�?k��y���jE�c�]T��sկ�����n1���2ౣ��x��2k>�L_A�|F͕#��p�֥���H#�%*��Sow#���H+�P����-���v5�o]{Їe]Θ]LD��<�=v���O�j!%��*���q��,±P���9έ�N-�Nf�9�]�i��������^�O�˅�'�Q�`d�	#��t�q&@�Ƌ�?�6��b���(/3\b�����-5y�;g�*���JvXB�Q��b��)���g5�H 1b����˟}�^�z��)D4���
��n7�>S��F�6��8'X�?���>�a���Y'd7Q�Jg�u�p[�D�P������n[c�F�jL.��2�#d"�v�j� �`��i��O#XB@w���n8��� 'v��\�e��
�r�i\�ۛI11��ښ�tg߂-�2��ː9Z,��.�l��܆�N'$�M�X֤�c���}�Q��@�4Jl��3�	Ƹ�rg.b�x��_���=�­r��R�7�#�I!�HiX��&�4M�=���Pl8T���y:��8$��_	��ԑ��T���9�O�8a��K��T]#|��'סk �����*�s��v9w� ��{�7ND�TuD��ނ�X�%�?'>�����Cч��!V��FI��?zR"?�N[;�ss(
H��\_��b���ᲾV%;,�4�t���P�L�[P_}Wa����%�X���p\Q������ ���b�*b<��.�m�D���g��� �_�)����دŹ|*P�E�?q�k�Q�s������~���}D��]귵�}�^��>�q���$/�9R�9=g�]���y2��j�9v��2�i�k�-��HlCv�ԁfB{�fK��AGX��ר�ς����׭D��/��o���D��k�%��-�nn.혟y̒�TlM�{8�+K�0|�E��ӟ1'<ua�Q���:T����w�w�$�	&pS¡��Zi��xf:G���+��
��������Ӹe�`C0.��b;�!<�) �c�(y���ʳB~>�댂w���6b�F�80xmV��a����8@5^�m:�mMEiX������2��A�m��d�NĮV��>�ri?sz4�3Fj���wK�$����<e)"È���a��#q�Wj�̦[� |+#��@ˡ�[��g7G��X�LI@���R�����N��Z��|#l1�fF�����Ze�����0M��@�p�&_=�a7��"h2�%�"����� <�*]�?�@�$G,Y]R1�׉�5ʟ�A���tc�Æ$n^�uq��$�)N�����9�tA�엖�4�ī?�5����P��o����<�F����=s�SN?l�4����
�[�GW���R����G_���p�Y�!���/Xt�V�f��Э3J���S�*O�mXX3�L ���Db��4�VfS7Hu,�s�6s�o�bq�H#�T�H�I���L���78������;���y*1#����+�?:@ߨ��րye���Q8�BZ�o9��>E�-/&{���&k�KO6	c��P%�=@�e�h���2=��s��9�DH�õ��i�Fw�!Ok`Hs���@����1��j�fz�~�o�nd�4�̘����Zz�c����:8�`=��X�E����j������V�Smӱnή�ܵ�I=&8�˙�]�[�]�K��\���Q.L`��۱��^ᝡ����o��O6SLWU�u#2�)�Gr@%�FrJ�uP8ډ-z�1+AQ��d#e�aL?+�4���./�]�a����Tӷ-F.)����r�e�+ͺIh�!�� �w���ld�0<���CQ�H:��n�V*;U 8I�6����}��)4z�cns�����Yd�X^qdN~+���F�0�9���"�`ǹ�*�+�5m]}��Κ�?B���`r�/���Ȉ��n8���g�u�dè����r	0-����ĸ`�3͵�Y2�Tuꢂ �*~8�j��kmI��u�-?V�V;b[6%�"l�ru\RT ��l��ۥ�?�c��{o�)��Ñd�L�u� ��Jf�Q����G�x3�Ξ��n��3]'�l%zZ�����z�I%f�l�8��}:U��ev�+4��%tS�ӡ$�����a;��[ÅZ)�3�����:���,�]�
J���<�%�cjd�/qW총�t��"/EQY[�v� 3�m�G��W]#s��v�%�MɃ-�0���%6�0K�*����ᾄ��a����*T	a�CJ)��W;���������2Z��.�a���8'��~�'E�_/�+з��?�a)x?�X���#T��	����/�m�L�P������I����"�X�۝�wkQ/	��;y���Jޒ8�F�f�ܣ5�H�֛������3�V#I�B
S?$�>m}d~���+����@u�ڛ�x������D-����4����h��x�KȤ�ׄdת��S�;%�ݚ�d�[��u�&��H���7�����b���yf$D�vE��j���<�j�|}�ҜB���g�󿏌�a�|
ꢒ ;��C��$�j�Uq��t8橄�=�6輵�g���V��]%�"j��A���?W��^����"mlC���`����,���,=�)�$I�����~s;P.1!�E�z}d��A��>�J�H��o���%Aٲ�`)%��"!)��<XH�K�^>��)/�$T����Ltp��U,C蛄��턬���D`����S�_`����9Gy�'F:ʕ�q�2���ӆɇ�4�<��F��ư�Z��8"0�e�!��R���U�N����u��u�޳�F�^N�z��eK}���1��4~}�)\�9\�-a�R�J"��i � f_O�{����8��c0K%Q��W������J4#�-y���1��gnpZ+���"姎r�gk$6���Z�p'(��������/��:!B���/k9e~��MY-'$Z�����W�7%4^s�r-<�Eo�⻰�oBi#����XXu��I6d�߰�1DPD �#��6i�8�4��S��#v���s'1N��
�g�!�/����Yβ�hL͓885鸴�:�~x=�$� �P�����[qWZ#�l5K֯���xj+i��*�]���xVC:z���WT$Q�`b�}F\mSg�_�ڸ�3���B�q5��&�6��1l��o8W�^<Z��F�O׹������xa�W��49S����UgK��rW�����E�=~��)�@)��1J$��N���F�-�D�fHqrFR�t�c_���g.='�>�N�S�o�#pkR���s@;'����d��u����^ ��:[j-��{�6��P:pК&����k�\R޶7ŝE��U��t;f�j�>��Ob�N˂��=E��y�g���',��0��M�#�Z�h�#6gl� T�:�5�������B\�v���=p�~oG`M�	�=,Y����B��ov���rϱ?e5� �_L�ܕ�F̎P��`D�05���J��[�	.�T��"v��c��J�� TƓ�?�k��N��r�-���F��PgNԡYj�C@��A~�3T
H�P����iz�o�M�~I����
X�iS�����x�p��Y b�L({f-��T��~���R��RC̚�kL�/��m����b���;�?����Κ�N�癤aT ��B9��T}��H�/.}���6��5���9vL�	�ή'���v�9U{bjO(�1Z�\���腐|��Sz��t-O�y�=JT�*	���O���5���,�l��aO.`�'�|c��n�_���$��!����6�x	6�	�U��ɿf鉜V�eab��r��C�!>��wB/�"縴<`?D���s�~Tp�(��^~��a��n�pGS����v�dN�%m�W���0����qBS5 �Bs�W��E�Y�1����v�K�r#���x��M.C�8a� ���A�ܡW�0���Y�܏�	��`yu_Ϯߞ�-w���(Ī(42P2k���*CӤ���`���TϠ�x7�[Tg��P�K�*�9,xF:���n]�����Ӿ�HoC�9��+Pa��Z:�}u#�	vN�蓕�3,Wڏ*�!O)�o?��Eg��2�
o��`H�I�~Uk��PgpC�¼ܩ��0Z|��<�K:9���f����P��5��;y�i�Du��`�3��xK�����<d��M��D	v�����Am�����2G�:�����LE��{n��i���mB	T����ϵm�:�5��#��L	(0)j��O=Q�H� G]R��s04P��M"l�X<>m{	����|�t^X-�'~t
k4�<�R���+N ���R��B�뷄�3(h�-��PW�[7M	����[zR]# �m�ѡ��\�M��{����
�R��J��^������}��c�V�R����9��tY�[4}��ۻ��b�'�$�z4��Yqs�7��n�v��sbn��b5�$4P7���S�z���=��/�EW%�wϝ!lrM���n�\x�(��X՗�=w��ʖ�6#���,��z$�K��}*�d*t' ���A����Gp�c�2B��Õ7�Ol��Po�Nl��U�7���9}6�����o��w+���Q�GAؚ�tQ�*�GWM����>�5s��K�O lp��S�{��2 Mi�#�E5��&0P|\�%�Âֺ��fqj�>��/�o�8�,���ݓ*�&m�����J]�W�D���߁�[��V�P�  ���e�+�.�$��bT�Cֽ ��+3�S/�{g�.f�_�¸���f� j�3'U2�Q��� ���]$R&\�<�X�1�:�$�	\���;{֗.�]�u{T-=�O�۔��T9�.�_�b!`�
T$��g{�쫦X��1��vL��D%]U�Sn���B��������-&�x�
��5�9hn}�F�@��s$�@�B��s%�����梵F4�8B~E�f+�s3��jH>��C���q7bՍz��G�0�|���<6�g,���� �+�v��ZN�*ٯ疯��@$!�����Y��Do[��
QJo�P�����ɍ�G�2�	+;s��5
 ��,~�%�t`H�#���y�Q]J��D`�]hPpy6�����sm���}��yv
��u��54�7��h�8X��P��+��>�W7M �867�E��@A�E��VJ�FN��(e���R�B�؆�4	'u΂:�3�X1}�}fA9�D�h8A�[7�HOv/����lRT7W�G2�qN;���\<�3=嘈d\ôzb;� Q�o����Sx!�($Y�u�8��d��E��U�@@Ϳ�,O l���8} ��vS�%�B�8�����z~�e���i�54�'�8奒f�}v-�H�*��ˑ�/�9C]�2�{X2�aQ6U�u�������ݏ+�D�����L&r���e�pm@X~Q�̪���0������鹣�N��'�z	�0�pI�kK9�%�+�|�!K�U`-�� �{!zN���.�!g(v�!,���'����~�q9�ũ1m/CAi���,� �Ӱ��w����49��s�MU���g�:0�j�ȣ|�ޤ֬lNv=q�]�c]��P:+��U�C0/�נ�\����s䓭(����+�k���홚�b~,�p6�N}��*+W%hp8#(����/;�=���}#t��}j@Z%J�x1#�4��#F����we�0��`�\������'D芨��5�|/�Ut�Q��~
lR0z+-/7�RziH���Ԃ�h�}���#�G�lK���@tz3�Ҝڔ�[�-s	eԹ��U��#?:�q���uA	�3��&e��Qb��R���Ǭ�]�۽��c2=&���,��tj�(���lfə��=ƥ�J�*$�^¡Jѣ2���	�(���}�.�e��S �߮�q�F�~�G�"��V� c1�gtܬ��I�vP3����z��=���z�o��&�Z��Y�fI�z�~a�۳���.آ��� ���/֒�����\H/Z�Փ��jIZb�"N�ya���ټQɧ�l�RA6'���>;Di��^��jV��U7IK���&�1�b�-|k&@z�0;��]�����hyz_��T+l��@�z�T�V�.o_�pc.�f�_��x�#�H$t��.Ur�=�ѝ'd��?��"%Ӂ�P��w:jO�st������b_��X)h�:&�h�3 }��������8NŪ4v���c��f��Gx��$o��xX���:�5�#0��/5��\[˹����Q]��]&hƔ�,�̥0���i�Gp/��e�C"O��dm�Udf���������]���:K��ݘ��m�<����������R�� <�T��1��|A��S ����A��RF �Y���%�M��s��Ա�\��0]6J�ȻѨD"�]�L����%^����ٯ��MV�����a"I`�&�Z6pT�t���>hb|�j��k�[Q#�_DO�w-�/�T��W���8�*�A�Xݞ��Dq���I;�^��M�;L�H�*����4IP�p�w��h�#�y�YԢ�;��N+@�Vӌ��Rѐ�mЕ�����@�U��޼ƭ�qo/�[A��s|��]�𭬽b�l��"*�0�߷��#%��e+�
���c֙���O��6=��g=����Q%��©8)��
^�s2䗳½'�$Nk86uDU[q��]�2ѩ���Y� �2��4]Z�N��z�oM�8�Ǽ?{�q]�z�b�r�l�qP�|z-P��	� sK<\{o�5����p��[w6X?���Z���8{���c��p���!7��(b-��2V��u�ݒ�>�T#N��g�3� ��B���o�>ցF� �|I[��<���ϰ�R�E����+��B�b��޹z��QZ�E�w��2;���A>�ƲtJ�&*���#ݍh���J;�� ���|��D_�Z���<�CA�.�׌�y��H��I�r�Fք��!w���/�]��zN������N)g������S�R��c(RyǨ��兀u3H*��Hez�~� @'�I�i_�#�ϧQ	!��x���U��2�A���e�s�I�voA��������v)��Y������֧��) =�y���i�fC>u�'��RWG@C������&��r�FT�G�v�H������6��eJ{�ɢ
�]�W�D�8��>�'���ƷBfg�p�(fR�R��1h��n�w���*U�aм��<XE@4�@U���woJ��v�>��(���t���*�{O�vw��*��:��XS2����̺��X匛����C��h�B��d�G�IkB��#�^  j ��ɳ��)��M�_�qj+Sxq�+��P:#���)�׌x���jhyV�^q�ޅ'_�j9�N��^��S��2A�����yvm� Hv+���$̼y����Bm���"�#�88��u^D}�F��^��- ���s�1큤��8ɋ�p��B�\��n�
���Ci���ZFt9�Te����h'�akO��]�{��N���*iH��|�M��R����Ro�ӭ�B��� jsJ�|�Mv<ơ���8d�V3�˜*��#jM|�
�;V�~�%�D��U��5���z�fR��̡��s�.C����8o^�IG:�ɩ��jψ(�R��of�#F�.%-������� �ģ#^��l�F�F���x��@_Y�(�$�GLo&u�g����<R�s	�FA	�~����t��uΦ��=nRe2�v��ѱBY�?�����{�������d~/��s�o�-I+�mRs���(-s>~�t�VT�<6�����˰ͺ�I;l�[��E/^{�&�� ���v��*_�p�ojWl y���_�bhc�W����$q�����%��c��XB�Q؍��v
��QWd���h�}=�p #R���b��]� Q���u��s�JG�ᔉv�xfI�0@��R�IҌ���B�,�#� ����_X�C5��
_a�tC�:!��Ձ����"�YS�f���	��l}�%x�Q���u�A���ӣ�Fo�Z�#���C�L~�	��O!'d`E����:w�$j|�h�.{�Z[]x��B��T���_6��=��ǈ��-��=}L� ��+O�<��Z,�=0v-��ꤽ�ir��=5��T��͖=ҋ�~^U�]�J�3�������Z�<���l#ec�]M��^T�:&�a��4���$A�~����6M沾ȡx3��d V%�1%���j��Gm���>6I���v{� ��uS]�S�6�N�I0��d���ȇ��Q���7�?�	V�4	b��5��p����c�mѪ��o�\�m�;���#����)�ze����
�~)���O�Zt��5 ''����|�y��q@x���&B�P!x}Y�WG�9�C�^����{��/`�d�I�kKx�Pk�sa"i�a��Z�w�qv�|JGd�Uג�(����S�ȡ������p�ϸ�*T�l�7+B�CK*�JI#�s�*�[���`@1f�Y<���Rl�2J/6^��FĶ��WA��#��n�!�᫐�n�
�)�GS��6N��iQдt!���F#a^�'��@�x�h�*'H�j�O������{�84ܢC� ~���#2q�<������G�CLc4�����e{-+8���^�xο�]x�� �l�Ҵ6���az�辦�����nU��AFX�[]%��[,u*拝�m*�T�+8y�c8%��┏��xe��wʱ���<�v�+hfe�c붇֑O��������eH6a�Q� �r�X۞��Yj�VT��H��z��vs�<ƨoPQ��{�E#%���+)��/k���(L�] ��k�XI��Q5]��`��y�P��ƥ��q� �?���VG��>z�E���}��T�\��U=g����>:e����R��/�I.�2����?�?���V�w&�yķ�>{�鴝�{�$�FD��j���y`re�����GS$K��� kJc�T��j�i(#$v1Pn�Z9�L���d�f�|�=g��J�9�U���\�bB\�<5���0Z*�˭r[r�j]6R<��:66��Z3:��q��x ��+S��zLȨ���4���١��V`aސ�+�u���k��tP�,�|ttM��z�:�Rc {�1�+�� ��@�"��w�a�Ӣ�lR�ϧ%�j`Ѐ�����[t�@�\�22@֝�_Y"��w���>�`��l��Vx���}�`���Sr�!�98.Y����R����a�Y�/�Ab���~�4a&������%�PX����edqJ�aw&J5�cpR(
F�P0y�Y��m���/3BD�i@��YthS���É�F3ǋ��ǿЈ s�=�om�Cg����i�w07=�]��<\�31ߐ�͊���G9�xb� ���F{Z�[����������CtXB��B)	�x��|^�1���l}6�QQ<����� �&��S����6���ʟ��oX�r�mT4t&�*܊e�W�lWiNy �ϙ߮��a+�i��s��`gCep�Iġ�N5���n�N���=Eܢ|�����Q���/����}E�{ϙꚔ3�_dM\��U���&�u���}m.� �.�s|į��1$��[cF g���׉[#��FT�� �ė�['W v���{N�6�X�8�	�Wo?�@��X�'�M+��-H(���t��⁎�K�ٖhK�ԓ�n�>�F�k�h���C|��;� 2
ko��v�]��Md�ê.�O`��|T?�l�q���
��� T��|������W+3QǵMq��>ʊܧ��.Wbҽ`;kYfy���=L��dGj��F��p��a�'֯Y䇗��A�@s?�� Q��u��1�U�rg���#�h_Ko�$;�,^؈R�E�7��a��k)��_�)���
���Xu�q�բ�2e]ߺ�K�
c�����Yj'F,.��ʲV:,�HUOЦi�����a%���|��w����+�O��jD�b���ջ�#JC��zK�������Y�1�s�r���-.�����"Ĕk�"�����$kNއy��|��Q�G��}}=��C��6�"{on`1�i�$��-�S n�G#�E���hF}������\�!|_G�k0aUF@�P���8p��V�3�'�.v�O�X���O��<Aͫk�D�;$���%�Ӱ;�`����KfR'��-��Ś���P���p�=Ŀ��,��I�?��MX����h�7*�AX0����A�Cb�0R��^��U:��b���I�h�-W�̕��08���-���E|V4���TCR]�t�����H��)����@���I|�.҉fu>~�HI �F�����A���P�9-\��O����p��~�K$����q+���5�g(�a�$V1f���g3r��f����.�sua� ��N�z�6{*��@Y�;=��$�J 0�F#L6iY����|"���޳�n��̳X����T���F�O�(��I�T�d0i>r9��C�=d/k�Np�S�Um9�X#�FC�G�)�����z���i�9�x�	#�A;+)��&�����7�X�nV��뫷���ʺ�N��v�f9�H�gs���R5)]�#[SFS	 r�I�?雗��)����hT%y0�7<�t1���8rUmJ
H�w�ˠc�xb�I�l&���.�3[~�k��eaC���h|ʳz���2H�ʐM����+S�t<O�=�5��>�5u����\���[dƉW$-T��ky]��������߹��&�ve��@ș8b�4���Z�S]�E����.��&�c��vι��U��}�k�h�A��_�5�{���Y�Qn��J��˰�c����DC�l��n8�z{�5�#�fc�����=���c7��@�d&��9<kJН�������2F��	�z��5�wU{�!���C=+h1	햪v���L�%P^:���9ㅠ��u[�2�p$:�r��oS9T�	J����B�i8H�e3�X��V+�^5�˦Z'������w^
D��MA�f+98kY��T@�)S����˯�{�ȒGsB3�k5����Y��&���gE��No.=[�Ƈ��Y�]�(F\P~6��3{mH��/G9�R�g�P�z���n�ea��&�V��x�)GO�+t�ۋ)_��G���� |,l��9і��1y$Y��m�^�ǆ@���,7E�V����I����M���U>�;���(ej��݁��Qͬ��H�ּ�9�^�U4�������gF�X��ە��9��ae����ǩ@(�^4z�Eh��Hc�z톂�S�t��j���by_�!C� NT�¨��YwJn0��;`� Ө=�W�4�;�i�����$���8y�^Yv�o���I��?�dߡ*�Az���� [�"b=�:�ڍ����$�����T�xZ�Z�c&�A{GF�c��aC��&�(��*Wv��������{p�5�M��R@@z�{�O��w�E��a�H4�g�"v��Ӻ�=��J���M���.���u�rQϼ�s4��}�N��ƠT
��,X4��Nv�[7e���g� 
ń���?��'}���7}��K�A���Q��v^TA^i�&q��&<eN~h��Ŋ�t�*�{�*��N��\���R��8�xi��S�S0z���[�,@~�0=܉�0;�G�@{��&D����V q����%{���)�Mj���c�^��RLR��pm���椄ئ���Ŧ�Ĺ���	]c�����!\�a���V�=�a�{�g�I��E��j��1��aꔗ(es�ꃖ������Ë*����1���V��2�u�n�����{�ۇ�K�Q��n�����L�Q?oP�a�$�ӻH��;�W�vݹD�B�?}����n:�rX�](Y�y_1o;�|:���!�Z�y��� ?ܰq{��e4�Ul_�N�k�̈́�-/�b�h�FBfoؖM�Ƌ,]۱Ay�,�~+`���xN_讑:_d��r���2�������ѱ�D�l��[�3d��
H�Q�U|G� ��<����MwA��5O;F��Su2:���{0�~c6/!��ʂ�((<�W�c��:�5�����K���}�u�J�r|ys�Ȥ_r����a@�QM�AT:Wֲ$W�"�iƅm	���:�N&�'���.�G�k|V �$�
���24<�1��h��88�=w�7y㷌a��&�X}��.�Η[ �� E-,GK����4U �2�:����X��%N�@{T�i�2ۢ�f���WP�T7	~����9��]�B�ׄ|/�KݞN�pwM)���՚��X�k��� ���uWAZ3�����t���rA�% �ԗ���B��d_���&��s�_���*��6�ir��D��p3�iYj&��Q�ͭ*qظ�l���L��c�'��/1�ա]]������-։��vّp>�vG^����+�:��F)Zi�����kr�4��nY%덕��%��-&ӈ�kG^T�}��m��,9u�9���-�ŗF��)�f~u��$r�VA+Zp����2�B�� ��ч��q�J��4��+G���������X�gR�K6Չ9:��8jT2a<e����n%Lͱ����:�w�.���r(\��g�=��9�!֢%�F����6�P]Mh�`�?����L�|����Ý�`�ȌM�6&��|P�{7�>�v�n�{��V����J)���Y�K7G�z^��˖}�6�����'�Zh��cH}I�vd`x .I�,Il��C��jGcR�1���va�?��r�jDA��tЎp�� �����?��Wd��[����#�h��eX7��U9A7"�09��d�������Ty�_84�oy=�6&+�s\��I�eB�g)@Vkڟ]�b*��L����_��O�qՊ��J<m��OO8��������{�@=�ujO�,������d M<y����vp��i��3##�0���d�1q��=�}(��?4󾀴�Q�g�k�#8s�,�K�{ _�`�B�Ȫ6�F]�ԙqo߻�1� �C��+R�ǚ.no/g��- �M�}h.��HLי���W��^��@��*�#c�Z��ڍ���6����ܼ�M������A��	�{������=�&\u�,BD'mZSվ"��H�����ouU+.��
�\]�Q�5!`R��d�zi��?q_S.�$n\�R?�X��H�4�o��do�U5���D�;ʔ!s��=ب���~�X�-��=@�c�K�z��N�iz���k�"F�gp�v��	g2$����O���Ǫh#��v�Ik�npiAq��N(-�!yt��YB�1�'�Ҏ������>��n����"kœ�Ub4��b�9M�����3�VM�d?A�q~ȝ�������~~E��e7�{'J��[��c��"�(Xۣ�%fiQ�"�}+��$�\B`��Tz뮂؂���C ��}] )ITt�xn�T^�8F�o�d���gVF8��[�X.�0�����%�D�;yM���#\�@ P������a��{���*�֯pF'��0R�dZ��(˩���G��V��r�a��:2w�y��4_^�+qe��F/��ˑ�Z�/�m�[���ÏD�#�2�]�eJb�|���	m
�/Zu��]8��VȆf�B�<	^}�C7n�u��7�����N���	����>~`�͓�|3E=�`�&����M�����B��Vːmk�$;��ɤ%��n����s1{�I2}@c�|�кx�d� ْ�:�n'�&�Hy�Nn���+�ZC�.��aA<0b��~�}�8��o�M8����F�p�?��^��)j��!�13���+���XNg��M�"��ʕX
{s�o�V D*�ҷ���n�&_�������Hx7apm|�?beU��CW&���/��u�ן��k�LWv.݀���}T8�3	*�W���w�XML�1%n��oY���j����"T>�(3\z������
h�j��c��d[��lŬ�$��ѯ4-!��}�~�dogc�}�
*�l_SRtJ(�B&�8s�'t+8���~���o8����cx$n��#�^M~�]7���aF#�6=^#�w�.n���w�})�j
Ϥ���L�6���V��;"���g�6g+��%�?~#�Y�(\���+���z��J�����pg��9sS1$?Q;�}���uf�J%��ϓ�A6�HK�'Yʇ^ֶ��5oP�����)GA
���9���1��u����"���p�>�Ԏ�-=�ä�n2��H� ��[��q0&�'{��9�ua$k��������(��<��JN���R���A������ ,UrZ8�[��>�_��K�`���ݲ�.��LZ��KLh���p1��Edr%��LS����W#�"�a	���ڧ�^��T �m�L6��xw�Z����55fP�m���VE��`ow�"`s�֖.\�lED���T#y�0!�P>ƥ����	�Sn�R?�2G�DLt�!a�4�E�vVןγ�$�55p��k`��_@�Ҍ�nl��d�;y��IWu�`�lB�\ ]"?��`0�u��B+���	۩�!bW��2��;/������Z�z��v�c��.D�nڶK��O5�@j�+��n�6�3�y^�>	��#5��
�7�*����ǹeplƶ��#�B�s�"�S"�Y� C06�;/�j*{<���Q���R/$����S8����:I)�T!�^-Mc��3=|�}_��F���Y�B�����zu��֌����1D�캮�O$A��5�A�}��f2G/n�Gma�8e(®��q���
˳�$?���X���َ	nO�kv3�r�2��зŅ�ف�4��mW���^���.��O�yl�G�E -���@����^bW$Q%�x#w�#���=�u�+d ��c�r���2b�F����_��q�AKީ�ک�	�Pr^��\Ĺ��k'�P��Î{O�5�����O*ד%�yyv�Е�e����&��]8�x�娛��}�Z���5%'f�V=i�з���#�f�9Vs��0�Z�-��>~�ȹ5�[��	�t�W����5��ov�w�5A��p��Jg�i��1�\ao���.��B1'��;�>]=U���[8�E���-�oؓ
ҴK��V��{�k�[�S��Lt�
y��g\�,G#r�^D�����ͥ�2�O��o>v~��݈�V7$���nX�Y���*���Jy���fR���ƚ-"���2]J:���Goq�L'�Dhb����ó�P�P���ύ�c�Ί���3M�S�ۧ���W������5vJ��2!�D:��Zz���6d	0���_ �,���$�}+���A������k���`��n�hF;���z��c�����5�C7{��,����V�`�`�)��I��=b���~��0��Ձn�W�������=��4D4*�`��:`�t~�B��B8-��¨`�P�趘E���b�
��)���g��	Y����p�s[F����eX�M����xLgO%&߽�q��4c��3��a%j}�r���h΢13҂�Xb���W������꟮���x��ǀc��qR�Wddډ{��G�D?��W�T;�#�m��:��6�8�T,BB�	�����7�+�%%2^Do�������dx@5��)ǟ	�7CA�/uד� �
�_�?+fu4Y4�R��w -U�u8�3p� ��5�BNJs׹�T�۰3\y����L������H�%<�&D�e��̚Hg�.����n���r��q:� k�\6���h�'j-Eݴ翷F��ًǄq���qމ)���R����1���⾭FC6;��3�ư^3g��J�ABH��ǉ�zQ�������L����y������=�Ք��w�%7��H����cH�`� �S}�)%����0��ۡH�
�4C���
�!���;t{���Nd+��������Y��tZ�	UQT۴�{u�`��
�t��n�c,�O7&�跚�ۑ�����o$l��/����QoMD	Xy��H��b��t���VS�9��=Ղd9��qYh23�X31ԡ��cyI����Z��J-�P�t������aj�x�%�����X$�X��
��HE@�݆0���@L�6�'�A�����Q��u�W����k�����el.>)6�T[6�t�P��(t5��x�q���i��ʍ���ɵW��2 �gRW<m���D�ӊ����F�}W�k�q�l5����p��_#����5�Һ��2��Q��k�(�DA˺�xiD]��ֵH�u��K�`dLH��O�� ��8��b�y�)� KI��^7(�&ӱ/i�f�+N7>���o��uGC���AXH���k�m ƭ��l[m����|��F�)�<�dd1�J�k}:����������!*5���c!��*يn/X]&.��g��[�A�^��)�w��4��ј>1�J��fn�t��� ,'���F��ԫ\0 ���XBͥ��o�*'�h� ��^\p��g ��
�#ׄW��5���^����n��7��P��Z��F}m�1(��g�bk�%����?MX�+�X��h?䄭��J�Wc{�h[._e���,5O�c3����$[�<S�ڹj١; �@$�%�+��X���㣡���IJOC�O��=���a�>Ǆ(L�U�����?q�����7�@
����ZESk��@�*J��DIu���ω�)S�}���I�j�2I~�?���t�s�,�r�/�@�̷��m�I:���G�d�&�1�gŬ勑�����v�-:��
���b��i	⌃ׇ��v��5��): 龰���N�2~��$ U��@����|���B��O�Oe�����qZ�����r6�hYA�>D�!�߉}k �X5��e���e�nZ���`�3av{Z��[�12P�f��6���_ͱ۞��V�n�E���o(L\���Mc<"h���l'S�h8����X^��"n�j�N�N��_���e����H���$M��(�}]y��ɉ��ǀ@��̑UhX^"ؤ�j��:�K6ƪo?O�G�l�3����;D��٧��sn���������J�� ��[bc��SЅπ��"s%U��Y����;l�u{x�L���=Q/�}U���}V��P�d8��ޖ��B�d�g� �������6��E�q}���GE���D�|����wG�61#�;^JtH��7,X?��Ts�|"Y។>uX�_����x6oq.8��蓳�R��ktd�gwc^����(,��K�c1�O�(��縒�P1�M�sRH4m;�[q�����-3M�0 W�$��	���C���Zj�2D�?�ZX?
y�9i9�E\�p���ew�t"�ee� ':mw�V|��Yv�V|^y�ih�|�xҚ(�����$I*��Ӧ���p�V0���s�͠� !����[��1��� �4��qH	4�G��
2�x�W��_>�l�8z�p�#tٽ}����ſ��|���u#�;�jh�M����8��eR3��!MȖx���2����S�'��_�3���'�ɚ9*.T�U�B�]�q��&mŜu�cq�>�}�ly�eJ��#����s;ǣf��|v��Q}���� ����"2V�kTU�����(��¶�sc��{��:����f3h�?,�	�Z�k�{wU�l�
��,�U#�	�JB0'7*�G��g�vJ��ۑ���[�����輪��_ga�DaMx�g%S/��◗
r�v&�ʹjal
5���=oӼΖ��u���/��!b��5N:K��ȧ�JÂ���B�2/K廜�z�	�Y�����Vđ���=�&8<����M�bP`:�������.Z�
5�7'�q�D�$��AJ���I��CK�����ex���ГRS�~�0k��1��" �ZԮW3�Qyb?nz�Gy|[�rɮ*sވ�w��iy��<���
����Ju�mc%q���Ɠ,T�^y�G��T��,E�5?�Un�)L��-��5�o8D6��k��Qbdwt&H�	��9��Щ.L�P��ɕ�w�g�J��v��!}K� �2%�N9ϱ�4cjOx�4��{���~�L��Q��V��ǌ`���œ:�D�Ω�ϯ��)0/CF.�Q��rじ;K�����VuΤ���*P���<a�7�J��J^�y�fO�[��m"����e���k0_��^�"��<�Tׅ�PB�
1gVu�\�4��Lw�6��a;8i�r�X�@���aYσ���g`�@�e��[�!B��^�����9ox#��� F��_�eJ,�b|�-�ά�F""L�����G���*@����_����:�.�4�8�[L��2�v)�gm �&iϨ_g�ʊ�-���Oj���	��/�a�t���l�_ZH,�q�,��qq�������>�8u��-O'KU��]|t�d��yjsъ*��^I�,u��u��Bm��r3�uMξ��-	-8��ع�s܁s���j�m6)U��2ۆ�Fu�O���u�Q/��@r�Nӡ��W�k*�����H$�h��B4�^��_;(ڈ�/�\jn�o+�r���v��Z�����C~��R!wd�8C�����˩��S�s�L�)����m;sӾ�'ٷ7FS�e0�x�,LsGmD�&`Y�����m�D���+�;Pf�sC&�_3h(�%gj�O?��\Y�Y�r�v�6G	PD���1�n�dKj_|P���٭6j�l��o�`�0cEaL<�gӖT�D�?׻�HW�*E���tp$2ТR�I橝pi��;��Bn.)B������T���������pI�%�z�x�׸�D���W;[��e��v�q)&n��hXi���h��fQ
�)�UQ�s�!��K���-��d)Y�@�[����9V^���r�E5������ �5�ջ I����Z�8�
�@���s�L~F
����+�]��>���I@]闊 Ru	��d��ɻpH���s�)��vBq�{ �jE)1��ԇ�Y����Vv�?�Z��=��\�z�"t�o붺��ǀ
�$ǴH��E�*���;�dQ�%���U.6�4�f�h}�t|8W���E�@H��VԌ9�Y$�(�,��üo��Ш�����~Q|�OR�Դ!e�wc������O)y�u��܄��ng�0����xS�C��E�7)���.�}��d����Ȥ���e+�&�I���h��|p�ԕ&�uYu{XY8&��XGgFU�XV���'�%�`��zrG��+�x��o%��x��-����p�w�ǈBx�_�v�#Y�����C��n�fCU;�Z|��3^���w�W^y���ޡY���� X�̜�}ha�D�Q���;�F��T7;�s�
p���̗(g*�߸`g`��lY�>f]C� ��3�5�U ��C�̊�5*���S�����V�O\��|�eQe-͝��x������������3Ox���o��r���X�V�|����s�$�yMy
��-���{s�B�@��ϭ�:{w��������U�h�u�M�B�(o�QUUe�y�<k��!d�ǩ
�"�9��h���5�������I��n�[�qRr����'�&{������ܱ����ӽޓ��@�M9���Z�v�i��%�O�n��k��ͦf��Đ�j��v�
h����C(4]��ӶL}R%XNqW�2��?5�h�و�����(e�f�/t���NV���9�o0N�}�Qw�D���A`&;�;����۩��]_{����R����	���37!K�"=��7>�r�J�4(�ZQ�WnN��%���gq-�F�1#��?�����Y꠺낑j���M�bYn����ƈF�g���ь��׽��H���c�����uع���n�u���I�`��U�I}�
���2��x��j5n3��-�x�4:�}B����
K;ߌ,�q�G`�wO3�Ն���tktBÇ���?A���4�1��Q����� �b�a*�C�y��N������~8�qٝF�Q�s*b�"�%� �w	��Td�C���>����MX���ag�à��Ǧ��ƶK�L�p"�AN�Б���V��0��-�K���;a�Xʫ�	��|
�7f��h���5�!XY&���rt�-�RX�=�nde��	}��|�ZN���(�R���c�d�δ|�-��`]���謕�"�5�z<0� �q�M��(�h��ɕ���d�=�dz�^�B�*�s�4aZ�1�;^���#���-/\����6}_������N�2{��&������J��Ac�y�a�Tb�^��ŵy6�J��I����޳�d�N�'�j����L���t%��n�"�fވ�<�.l��&�ݮJ��N�=�q��ΑZ�p�Ƶ"�ݎx�U*��ϱ1�>�����T��u�zo:x��%J=nJ	e"���.>֨_Հ��3��e�Z*1j��F����y����ߧ��h]��d���sL'3���O>�b���QY�0��Ñ�p��������H)R/x&N�����*�G��!7d�b���[����+Wg��$f�w��AW���g���R���Cy��Ɔ�S�TC�����XVF�,l�2~f��ΰ!���D�p�˪p'_�L�~��������7���g�
�y��{k�>-.�D}h[����XF�������9�v!�D҃��Oc??7'Q�H��x������'S�e���y��3��Qެ-&�޻Y��˂�.�$:��|R{�Ё���v�$���V90\2gcf��XEM  J�(��Sc�<-�٬¾�u��X������V܅�*Kb�Q�Gt�p��s�zX���5��0Tª_��_��7�x
��]ҭKk�'���<�k�Du�}���W�ө�]�Z8m�m*���YÀX�Ր ?�L�ǀΎ�MT��������g~�o��^K#>�[��%-���1���'t����}���+z�E1O�1�Bû�5��ʃ�lEiЕҒ��x�l�,<�צ��Cc�ys���l��E9n��cS����sy�j� ��w��� ��]����j�r��1�>��`�d�mx���>[���"n�Y#RB�:���'
Ok�ݽeQ�n �x��(�#O`%r�x�3z�\�'K���K���t�+L]��M=V�m��=*sɛ����c{����-t�ߖo�͓�d�«�����Eq��a��.�ǳ��@����Ի..�Y�ɠ��I�U(x3�d�&Q��ϕ���=�'Z[5�����ֻI%g�ݗ���M�<�13�+��X�b�
%4�����:-���F��`�K9����8�\�M��]��U/����\~��2q��Po��T ��Bo��W�50&��ᯏ������/d�\�}��1&z5T%?G�����~���� ���0��-@��=�Q�wl>8�D���<���wf����?r���PC��@-��P]�E&�󳍴�9��>�e����Cw�C ����sp����&UXDb�$�R�#����	�n�x��,�g���C!��T��rݙ	���v\%�s\��{���>�Ak�.OҴڳG�Lg��a��+(�� �KK�L���v���h��]矏��Xq��Ԋ�ZXL��L�՚<S7��T�f+Z �om��
+��mL1)�#<��`)�
	/�0��$�ru�l07�?�;��`�,������*T�z6�k�e5��O����hR���E�a;�@�'���D�ut�M�����]�^����o��rD���d_����kJ��:�jì�	-L�	��g]��Tm�k.���cy`4���%��U�[��e���鳮	���gu[�^5�o�����������Hg���������e��ƅ��rY�p):쉦@�->B^H,|W*>L��-*�8g�Y����Dw�L�H�a(��Y����܁�TU�� ;a�5�p�&}��1x�f�q`M@�b�"ɰ˄M���G��8��*+]놪����$
}�@�3�}Fo,9� Wz�*�J� �/~�p�+4P�)�t�$ó�s|���[�I#���U3���� m/r��o>�iH�.
4�x8��:_-G�mAg2̼	S.�6�Q�E �.�iO�����Pp�q6�q��1LB�4�����q~t�fD���,qF:�aR���S�D����Y��JJ�t$JY��G�*A��;V���j_Y��=�N�	Y@$��/@��6��޾�|��y����2���,
��U����j�G�t} *D����P�vtW������|8�������EU��p4[��^��u� ��+�,N��
�yBQĀ/W�������9lO�X�d_�`�'�����ӑ��3��ǐ��*pj��/�%1A��́�Jp�m->�߀���O����t�?Nmޙ7������q�Be&s�/_6Z�s0!9]=���7��6��e̦��EO��/L��@�h��4�9����<E�M��"
.����s�)黑`BKn��.ȌT�m�LW�x���Y�e4���,L���)�1j横�ݚ�ۑ:�����ɾ�������w��ܩ���"X݁c��|�L�G�-;F,&�I�B�����~p�v�A�S�#{�x���)��y�^�_j��BKM!kBN�ǭX�&�Y�r�I���OP���r*��!/fI�67���@��5 �L�c�׹Ң��3�l�����9I�:�5��20����Nd2:A�)��Ճ*f�F	���پ\k97��g��5��)��>/\���Eތy�a�y��|���4�q�rkٵ�п<�^(�6�o��{>#������v�FT�o�8��K����!�>R!f^� �-|��7�XB/Ԕ�1��k����1�Y��N��K�6!vS�����5�ܾ9��t�\�y�M��oC�7��}����5�LV`��.��^����+|�h@�m�T�<��"��Iy���6��J��/�Z�-�ѧ���T�$p�	����� ��x�\^��UΏ�x��������������	JPՂ������� �SR����R�%�X��ᦍDЖ����|�񗝪i�r�.���%�y�4ĊavO�#���g�qN�Q����O:��kTSR�ȭ�n/��_�"Sۡ}�@Q��]�Wr����*x�� os��`7�U?���*�S;U`[�'Ɏ|S��I�*�!_HAe�@�V獝cv\�$'�����h��v'�d��8>�o�k-7}��_S?��<��mcc�:�������z��R�ZB�)�IIй:��s���F�!y�!ښy���[��vf��~�l��0��~�>Ѽ�*����p����RcSp�f��>��;��n�C�]��QWl��˫�= �*�&���6�i�G �UD�	��#�*K�����?&��\2��e1��+�ԍ});X`t�tP���<2����u���_ޣ�P�A:�'��61��I�`O��%��Q��a��Y��2pL���(��Ϡ,
��ڪ�%ƥG��2��!�TM������jt!�{+s;K��0���VNKB^�,b���.�I�ߍ��ۿ#��{w=�]d�<����|yH3M�*�hxEE�7�S��E���M׏h��.
��D4��:ܯ����Ԏ�}����&G&�Mj��x�#8����#X��z߯E�jQ�><)C���ʪRŋ���fk��i��]�X�݊�	S(�aq|���
Fs��{b�+@�a5���q�)���o��}�a�D�G��j�=�q���_��٣]�Yn���5�h� ԭZL�]r��5�Pe�м���c�T����7:��X�m]`้�<��9��b�E�i� �Li�ڞm�<���&�^L�3`
"��i��o�Ǥ������� |G�S����x�:�J��[�Ҕ�p�-t7P5�N`��P�.A"i5��ܫ��gC�����u�X�2��(p����)��Vj��r�~P���A�,�Y��R�>�dy}���%ڕ������Q(Rr�RV���t{{UT����%Г�K<!���5�~����C�n�t� "�6C:�>�M�[Hw��!G��jAe��>����K�4l~b*M���La�S ��z-�i�b3\*Y�B��0��
��4JqJDc�Ȕ��nOO��f{ا�.�}�m� %��o�A�D���E�)ף}z;ZM�Of!o�ܸm^�5��I��8�~����7!q����H[j��ܡz�]�M�?It���z������6�\~�Z1�H�

�QZ"{��w�ڋ���o����n4O�Ur�v��N%cípO��%�ȇ1����Bs�A��1�����<�8w:���Z�(�V�p��	ئ�O��?������T�=m��b��JO�I�]�	K������������I�tg'&�����`�)�h�������9Ԝ{�ll�{�nT)�8C~t��K$�x衑(cD����,s"�"�#;�v�I)��^�O�`�ʕfRQ����_�mV��ǯ/ǌ
�2�����tM��P�o���^�����\�G�{��9���̃�b�Y�u�v�U=Zg@�%d��gCI�Z��"�S�μ�l-�=��l^PN��?U��Ι\	+��X �"��n��\�j#='#a�N	3�5���֭%���-�I7����3���x�}u�U�����8�sC�)��(6-c�t][gk����/��
�b�kL��Q@���
d|�mV���5�R~�5E����!6 ��|`�iK�߸����-x=ȓF h�X'Ѣw��Qf����9�nȚ.����Rz��!��[��[	��,���a������0n*D����G��@!XG�ݡXy��u}��4�~�(ⲙ����V�d�ɟʮ���P�UtޫYc��(�z7��&�	�D����$��D���Dj�*ĝ3̘&�����e�[��n�ZN�͛E��z��"sl%(�4ET�ݱ{���'(�H�;"6�
�]���5�>=-��1����ڐ��(k�Wp��g3�z�c�$B�	!lE#m ԝ9x��R�m ��������v3K>�0���K"9陌����/�e�a��(����tJ^d�,O�V)y^������N�F�����k�%�[ sHJ�:�	'���J�V'XB��̀���p<428�P<'��A����rm��6��erʪ|��s�P��rgFWh�:�"y��D<Jt $��A�q���n�а�����#yRkKT����B��L�}���Es;x.�},?l]�n�%��j^H��(Q }�8�=�n�1�
|�ȌJ��`����pk�9^-C��4\䛭.}��VS��ж�����؟2���_6v��1���4�U�d���ȯ�6�^�o����̠�Z��"(z�֋��4Б	8���M-:�~��'Ԥz=ٰ�P���qE��I5AJ<9�� Q��(龴�ׇY(��D�_%g�kXl�9��X�Y��#�~ֲ��ú2�k:�K�k5.�(T�& C?⟴�������8��DTf������bd�"W\h�axV��TG�V�����:��4i�ES�M� ����@=�)0��XW�T�?E��V������ez��Ap�9"��~"�p�W�0���ꈞ�]��@o��
�̵�Ր8J�0�8�`�f�'kD��&H��;��֊($�]2�*�Hj�b�����4��Rq) qW/4�����X@�����,�'�H4r���]�\�F����F���&[y.�PH~{C:�y
���
���d�yTu��PaO/>w����zVc��P��S���*�|�#�
	��Z�ɇ��Q�7��H��2���8>�3�\z�$����	R�u�;��#�4��*�i����_�.�p�O4���xSQ{�'��qH��T��~�8�P����!G��/V��diB�.o��_ؙ;�[b�-!4�}��y������>�pe{l�3�:�6|���{7wrI��(�9 ��=����>������I����?Kg��?�"a���`W���Ul��&5��#t,�k�J�����;��7�B�#wKQ֣��{�lx/���x�$żRIGNM���F����|S�5��#�zw�� n�̉_ȱ3�*����c?&cAG2�'h,hh�8b�PT��O��2����VAЂ��c^��*�#�3�CH^S�ӱMPB��E2v����#��5�+�F���)�n���yo�LgH$w�r�ߎ4���-� r5%Bvꦻ��g*�*�B�e����;k�h{�>�(h��,"�Xa�ZؖD
֑p䡒v6��X�]/��F������6���1����X3AD�27���د��+����V�P�H�6Q��ap8�_?�k�{����wAC��t΃FL�%	���(���(��C��$3��'�
Y�� 4��?}� �>�K��R�R�ź�X譍$T).~k�jw�U��^|S���"h��_�$���H��x�Z��(�to�q�ڬD(�c��U��u r�cGMلOc��$�0�t@�Ҟ+�30��(7\ ��v%ǅ�C#�:f�:q���8sXS���R
B�`����C��V��q"�7Y�y�h"C�'6]��ً�����L}5���{m(���{�O�[rBr��'Rz��Vp�0O�0o�h�.�Y0*9��6���U].&�����FN��+f8+}��������dײ��,G႟�x�v�
��T�*=�`�z\����x
�rO���rͧ���U�w��
s��ם�~V�<5)}���Z*׳$ �hZ<+��źK%;7�tB�Ƃҹ�;Dү�;��,j9����e��R�w�n�}]�M;g�P6Is���pnT�փ��t�g�i}V�c��tL�F�+Yͪ ����.��C:����xe��;��˯�$��)���/;���y
FC�Z��-hÜ#͓b?ǔa:�g-쑾�VYfw�:��'ɴ�۠�*��!I!�J�cg��h,'��X�x�gD��)��m�A����N�'Jf��|�J�,}1w��z�#û�����<C�[j|K��'*�d,m����c��;A*���2@�/w�Y��
,�9�z��0l^�䄓`�h[^���֧������RʹJ�HK#���σ֩ą��"��!�?�]�[�+u�.z����C���+�����͉T=����<Б�7�F�9YI�ee,�6'P=��$�����&
�8����au���u7X+cDF@�H{�쿾P>I�uLA��[�zq7��ͨ*��,�!#�.ZY�QI����Ȇ����������x��b,�n`���5Ģ����-�Fzw.���������f �g�U@?U���yB�z�x[�N�S����Sq�L�J3�$+�;��P��Ό�oe���D��f��w��ѼF/1�Xw���}�c�~m��'��T�u����8�[P8�E��:��	-�a{w����Ҿ��xg��Ka���	`C?�rG�;
#lH��t�ۦ��T˖jS�H�w��?L�<��\���B � �Z!f�>��m\:��t�pu�_켨C�a[q�zJ�vuP�07��3G��JI��ECgCO��v̕<�z܇�L+���n�3N��j��R��AظA���xD{�ؔA�xD 9#0�n�~	�9s�Iz������t�.nvH2ba�r��Mu�P���& nn.�}@7�d��!�l銼	F!��,bQ�d ��
��!�gAe}f1�$\������4�R~�)��	����]��S�Pӈ'��YKIR'�D9j2j�mAA�ʌr��hyd�Cu��&G�p��*��8�V[2U�Y���F{�����Y=-G�6�k��Y�P�"�l�<^?A��Qx��H�	R|1��4S��i����o<g�@1腍<Td����󥮥�R����W�;�m����L�]V�5��C�1�F/B�ý�w��u`r/���Ν��Y�+��I��5\�{]8��|]|���Mk`-�r�J�,�i\�hǣ&�Jҿ9��:�;�J����jIx�@i>�*�.��%��=F�cN]�����]�)�X�|VG��i�yV��[j}E>M�� Е��k/";M��N�%��/@$���P��T�Ʉ�bo�%�N��k���%�u.��#��{�	qE��(��1�E�O(rE�'���5��) @C%���U�!�����:L�.jr�u��V��7�|���'ă�1��K3(�"�ZlT{!|ۑ�tݡ����WU��R ��F<�փ���ʼI�<(�{�Y5����yV*m�Qв���Y��dCc�zx�h��{i�r s��S
�1�r�I"%���CIan@3�����4(��:C�Ht�r�4)���J����2AH�D��:$�Vԣ���7�'�e�k��3�e"�^vk��1�\� 7�[�m�Ԅz.�������e�$��'9FK'�zo#���'6�w�����J����I�s�R7U|Q�*�D���d��`���)]�9m�UA��n�{5��-s�MJ��Yo;�*\���$�5��N[*kq�|_��2;)Շ��uۄ�ϫ��@1Q�,�=D���=y��wI|,a��7?���3d��=��5}�D���O
��}kd<&�l��M�J��E��0�Z�����W��e�j��e���?�0���1��	p��XuudH�vS��mX�iy�=AJ���D}���hfKIQ��ݍ��K*����m�ꭓ�.o�B��(��0'��i�Ѵ6�a�Ћ_U����ԟU9��~?|9��,�5.�,N��cxK&��R���J�E����~3'~��|�y��P���x� 71�=�u�?�V�H�!����C.̋�@�V!lo�(�j������6�Y0�Ǻ����c�0�$�~Do��k}`�z��{���X�����C/ؠؕ�&��������Ƀ�;��Uw�`�����<�݆#B�Ѻ�{�Q�l�K�&>�#K�P�q� =�?��|�� ��Q!zJ���ACQ�с��0p��2���Jm/�]Uqd��$��4i�w��,���������&��,^1���~Fб���$�@�00e��|�óU��Фj�?ѥ[��v?����魫ߠh�{I�
�LԾ��=��y:�`=���P���ȾUR��^�A`���Q�N�Խ2�4�����^��!�jv��f�|�UO~�m�����oy|(K�<~�*6NJ/�3�dv8ObeS!��r���D;���J�V���e���n�.����U�{?�v�R��!�P�y�j�".����5��Z�?�N���7z'������M\4=Ưr����ܼ�(�h�dT�]U$�DF�����:p0}8ū9���Uvt�i,w+�@x�8�8��n	������ĵ�%C�TV��#¥Zh���� �f&�ov�
�(�ρ�z@�����Ov��s��f�.B��[�B�k��x���!�U�#�]�&�ѳ`���J�X����OսS��;�o��p��}��dC�x	[?��9�(��&�1��G�yi��	l(�Qء���fv���U�F-�L��0���\=1&�C�����8��w��V��n߽\0��%v�$iH"2����ޗ��p�^@�e��Dzc�D�<$h�`�2r4W[�L�w����Л�X���z^d&��"psd�����ƨ�E�7mt��$8�!��lUQ����C� �QC�75A�U�Ƀ��� ��,��5��i^WH�@S�$����W2��������8��S�4�m{j�~o�:�#t�tb\�`tWldU�=@Fr#4����O�"z����)���z���h2bHl@Z7llhe�#RX4�ȣ������S��d��sJ���(�G��>F�Œ)�i)�SC�Q��k�W��!�Z ͜�lQ$�Fb2�>��><�N�G^u����s���Ì?�4�ԧ�\�7�����+�f��~�`E��~a�YmT�S}��2�u�8��Lk"Hv|wj�L"����[�{Z���C�54�i� �U�@v2��}[�DJpU[�U��8���Ԡ��0���m'�yx����A`��_H�T��"aN�����Ǵ��rxˏ�uN+����b�txbs!,-Zy	ܛ���U`v�ol�J����,t�#�I��u�k�B�HBwg�m+�8w�0u>���k�VHV��H|��26�K`�"�}�����-Q��~��}�Z&�	nK��
S�z�����|o���[���"�
��КYئ�G��i���{�1��9�UŌ��R�gs�q�q����D��U�zD^���}��jpnuB�2�6;�5wZ*Tr&�����rx{V���qO�+k~G�H����EK�^��dg��h7��vT�{/H���*N�K�($0)Jp$�ວ[�Կ��R� ���ze@��*вƹ��1�;6�t�G�m��2�5u0�6�� !|�hi ���[�n6�>���!lP�H���÷���-�Հ�_ĸ����W!r�[�5,T�J2>���zk���ݢ�\7E�@g��Ym�C�@D3�f�x�gv��Y䣿x����BM�M[�jvUֆZ�ď��%�}�bЅ��m�	��E~�ތ�{�Ĺ������\MgvQ`��-O�W�qϽ�t٧i��nO�n& $�('�Q���뀲X�:��h�`K��-��#��(w��Y"s}��Z)CJ,iY�;�]�>���fr*b@u�w�M���^+�Z��a7v&X���5�w�j���%<e�QG&�k�Y�%<O5�%�f��V��o���7��@c�yC�>�~2����Yp�h�|iQ,�L��'��Wv���S�K���n�W�7~�_PXx�5j<\�X�i�g��)���1�[�����l_?!N>yN�>ln�u##;��9��d���`�S`sf;tp�0ΐK �	��M��+s$��H��'��!4%M��pv�Uű��Kq�u���)�#RRJF'�uj�/����>pa{�qHՂ\i#�=Ҋ�/w�G��X��/d���e�\�/H{��
��Bd�Yvr�ɺӬ�ZK��X��f~�cF4���Ho16����������fk,QY�����ze��c�jB�/~�q8./M��j<�h�Un���|�\G%�w���y\�w�1�e�O���谆؛j�6��ƫ�{�aab-G-v��5�#tG��\�8�)�T.������P�4q7���!_{��o3�6Ͳ�2�7o�(�[ k4� �}� �+B<��t�V±ږW�Y�4Ht����?Yk �&K�\;��o�eU��i@�������co�BЂ��؞�<�FN+�S�Ae'��0�#_�(��6?��q�@ʳ�]m����ut��kI�J}n��j��c4Fp�����0w��a��2\�J�� ��V_Ȩ��X�]j6z�R�#��K%�`��R�?PXr��h'v[^��mX�Rl�)�jD�3u�P��
_Ju��]U��]M�@��:�:�A%�͏6�����4|1�F9�r���/�s����<Z�2J��fJ�����T����O�0�jgS34%�P���K�A�c?OC��z.��E͜�~��G�O�8���	�Q8�Ln��.�<�P�Og�7+i�f�	�g�zÚL�]f��z�$�ȇMP`��Ŗf�,r�-9V�UK2���xa<���ϻ�in��5�}v�?r��j��t�x����]�ײc0k�8��o����9+�R�(�vƐ��%|z�!5%8�tl���yۡ̓E���l��<����PSPlz�D��Ռ�¤%�0��fX�C28���^�Ꭶ����[���>�k��p�=��:5�a0>nB��<��L�miguS�Ҋi��b�P�X�����Ҝ.y��O])0��u�kд���*لoA���z�ԙ>�^'H�<��DAޟ{�Y�[�����|�p��4�Y~%��.\M(��u���m��c ĩ%��v����/jM��h���iN~c3����tЇ��ko��ꥯQz�7��S�L�?-/�)�8&2��P-[�y�F5#��\8k]��d��b>��αu��^>C��u���@ߘ�,���@C�52E)�4��}ffwC�
ӊ��D�����b��;�:��ᯔv���[O;(�����|͆�_�=Mfd�vM�c��D�-K@�VMzN��8� H}i�f�􉤨���T��D�Z2Š��ڨ��������7��V��+D[���T��u����-+R���G��ɿ�-�(�N:��
���hV훣^�3���)��]��5�u#5zL��2��>�M/��ڪ�@�|Q�#ת�`hN�z��U�n��0��cB'�P��o�$�8ӳְ�����u7�q��=Yn�*M��N͠��ne ��!��*��6+0�M����6j;���>�bg7\/�1�� ci�������u� �/2���6�7�ۼ��1��h̯�f�d6��S�����Ul�����@������\����q��i�Wh���e{� �����צ�� zW����ZޑE�j:�Ҭ"�[ج�����!�ypF��0��c���|�{��,��l�f�q3�̳_��ާӃj��ªgj�����;�;��i#rq�ݶq\'z�!:�8���}�3�#
{S��X�XnM�O�1�SG�<���x���~���@ų�wygp3�T8t,�Y�����f?'�	
G�Q���`�ֶ0Du#H���xj�xj�������uf^
U<b��1b��N���J̘�+��N,��d��|OX�WX�tu]f*õh�|�wm
؞W��N�����/�Qs_ n
�ɹ9�C�M;Yi�B�QŦ��;�b�B�#��tg͝�D����E��2��R
�z�Ҟ�-ն�R�1�ׯe���EX��G��`&r.��n��wpT���Ȭ�>�S�j�(k�mWc�M���a]O1[F��"z��Z�3�̥���M(��t���꼀hԐ�.�����S�i�V;K%e�������TZ*�G��U��B�2;��DE5�8���2
���LՎ|�t�jȀ�`b���a��%�9�dcͽ�ӊ�0��.4XI�����W��c��t?��(#�4S�{��3�r�l����ʻ�ZS�J�`�aLK�<���I+�4 �����%�L�]�R���N�p\VCKx|��'o�@:��e���,��5���i7��*m�NM��AoW*�A_�2KK�ŷO����v;P��V���	j�P���rR2F ����Gm�2G�҃=i2�.�xh�0�I��[�oCh��� ݍC�dp��RdXy��q+��� ���κ�E1�O{{��l�؅��rJ�+Mn��i���[z
cw�e!����	`��D�H�1��N�.�֙���<:7d��%e��~�潷�剺|ll[��ztǶ\���:��Q�@���Q��^�-̽�6i؟�N�����ud�a�I���3�
/�e m��w���Th:��e_�>{_K��ڱ"���.��7`Q�9�I���R����N�$5s�%S��p!E��t"/u��w����ȡ�<����Fӆ��Hb��8�q=u�ey�kPwz���g@�X�;W�.0�#T���~��oI��99̣�2z�S�1~�	i�+m�{�nm��˜w���(���������d\k���Qe���˄�Z�$b�Z^~�oE�[�Ʒ�0�t[�@^.^���ϑ�a����{3A�����:qH�K<ZƜ/et���O��dL[Ge��{Hs�Ge@
6�Dl��MT=����pE4;jd F�!�9��L�8�kG��-��&@�s�2��������֛��{I2����۰�\�d�YPz@8�%@��g�4ML�j9.����E����OO8#�N���ka<kp*���6�\ֳ��2l�I }Ϯ?��gI�.i�|l���f/w�~`��!w�$ҁ��^�	8���/�uzս�N�|�D(�]����C����y$�o�ov��x��,�^��6/gN�ت���?��ޝ�H^���V�A�
f�WV6��^q?CA.;�\��Q���`p��m |�e��K�-gP��� Y˹�US�gS�:j��/2��%P�#�D�8'���`Ṥa��y���"@)fKZw�ˤ�-fV�nE��d�e������=x5J��>Z{Y$��� 0d��|���;��NM@'� i"?�*�WRc��So���z�ڌw�l��/���\�g�ҫ��G����I创�
���G��d��C\��4��qך5�����]	�V4�"f�1���m��#���Cz���>N�]Y->C�@`�\%g{��|b����j�)��	ǼiK^�_-�\�P<5f)z�ʳ���?/C ���MG���g�����+;�޽�G�٭�C������O�l�i2�5	̫�n���EzDN����D��evZ �PkEx�&�+H��&M����-�~�7s2]�����ݴs�cug��Լ�6�z����D���G1>���"��4w3Ρ !��2��wԂ��LRM�����8�~y2��,�Zjp�諾"P�71���=E��g��uUr&j��6i �����O�@�Qi��rDb��p�	�w2�/�#�>�L�f^^�bħ$�AH���,�V@L�D�F�p]���afe��_r	>���Qcs]��cgU��`)KRC�S�_���[Ԋ�@]ծ3��@��+����K�#� ��XY�[d2ز*\g�y�������n@���n/'�+�u��̦�8m%=�K�ʑ�di0x*�H�!����Ҕ݀"DԆ�c$������_�^��n����T�93d@=Hl-	a�Z�t&iǴ���q�����)ox_#��vq��S�zF�p��:v�,(Xyw�c���Fjt���j�-m
毳ᘹ47�r�S�"F�#��'0�����~>�s�;����;�a�S��n���_�\@�n;�u�ཻ z���7P��P���*�m[�,�u?.r"/i�_�g����9�gtnƥ���D����1��ny���)��B3������0�}��h�:n�#J��e�T�m����6�{(Ǘ�9|�W
����Zn��X���TKV�;���ű^��G�a\�k,��b��5�Rl�kr���^�5�Tk_
<8� �j�W,B4�h�y_t��'���z!����ի#�f�O����2ڏ׍&zG3�,�7�s�l/!�E��d	�0�2��!5���>���iW�"l���X:_?�R"i�$��{�N��k�9ܵW\J�����k��+�(Z����b�*P~���������4��7�b�X�?���D:̲��0Eɔ�F�ܽ �D?.X)9�l���7�����T7���	�N&{�{�'�	����c�=��3�ղ��G���k��T�5�M�.¾�ZĴ��E&ݥ��1��ߌI�D2��|l���`{4K^:��Qd����菓oWŚ:���w���<�Ǵ��8�E�%�`��C��)�G�lw'J/z��
I����8����W��Zu3g:�OW?�w.�^��7X�V}����y�0S�2��-�d�s	��;��o v�9�{���T�H����nj"���B#0=T��-�J/�h���Q�C9
+L�*�}��|�W�8Ħ�b�w�E���	��h�d�tms�?b�?@:؊���l�\q]<��g�>lU��]��ϴ��y`̉���U�K{q�0���-/�����5f����q���Gi%��*6�o��i�`����i6�9��c@c����D�.���z1�bC�)%�#=��c~��s�C�X�?'��J�Uy�6��F�/?����L\L���-�~��Q)JxNiF�	ldMP�wqR�Z�*����a�s����_D��"����p��a��X{���O�YwrQ��Ϫ[���u,����C��-��dԜ, : �fE��l��Ka2���ze
�=���S�{?
�l7U��E8�V�d��E����$)\+�~�H��cc�V\b�0<%����HyX��|�ɩ�X=7�ڢ4
�A�	����$��)���9}Z�xU� #L�,��u�������鋊L����4���R��,K02�V��u�k���5t3���3��bY������j>�3�0S<��߯�}oz��J���6-B����O-�<��J)G���`h�UndQ�/��D��$���>���`\v��NN��d=�����FV�7�K���w��t���)�v��3l%B=���4�'��fK4���!����c_y�����ܐ[iL��Q�0�$���?�g�(�~����,��3d"Lk�x�%0�@YҊ�W�r����˘Ed���]">�}��+lq6�a�#�W�Ӊ�<R�-���n��;t��U��ҵ�oZ.iY�qZ�����T�!�e0���._��x֒�t,��t�K�R�W��=��%��^�,݈h~5+���ʼ'@��6�`ˣ�+?;�����S�)Ժ�Րwa}�9y�|��U߫����4H�w�#�v��*�yO>������6�Y���&Q�rj�8jB�ty+|�ىQ�}& ��@Oe�r���~x?ȵ�y�IC2�̢��@�8����`�6�8���o���[W�xZ��;�2���r��	G
��M�[c�W��l\OP���`�&�"z���P	��(����E�Io?Z���

b)��3ͻ=;���V���:^�	.�LD�5�L�ΐ����ZӞ�}�V[U�_����h�o�L�;f
'�O��pw����X{"����c�����\���H�z�DA��ۂ��`?���Y)�7�
�w?}-��R���YtM�(���9��Y��<�����E`ݜ��cr���j�#=G5l���H�
x�#��dK"��hAk��rn�V_[��ڇ�b}����8�a`5����o��w��?�p++���Fj�7!OA���:
+�+�T�"��>�N��'��Ez�dI��Bd��d6O�i=hT�9��cZ�/�*�&f�y�? �Z�	` �N�2�I��L��+b���C Y�6��J�xErqw���&�;�v^>���I?�z�~����F��*�� ���Z�Wu��Ē�3�Ɵ�ݫ5��v������\�v�@����F�J��v�&�σtTXT��~Ռ}��	<��D,,2S��'6�C|���������kv�y�Ŗ���x���o��>��7��-E�&^&�	�ﶆI���@HA�*q�j��of�؎�e�[�A,�3�����o�N�5�p̜�V`�7��I�c�H�5��>�b��)Ǧ�O'bLK�3tT��LE��]�i�DQ%A�'Sep>o����<�� �
���p��"�Qժ�^և����̅�h�'���0&��c�ȇ���Z�߀����<��ٲ�]h��3��}�HT�ӂ]�����H���!/x��w�'���A��ĥ�O�@>ș~[}�N�����F�����0N!ٳh4�p`%�E8����[U�3��[��aR�G���e��N�Pbnxu]Qp�{�DnV���S����ڬm8v��W��F�*�n��#����0�M�CB^�5���R�X�ę���j\\fD��t������V��"���zL
_�}����P�|�@X��8��������!!����~�W͊�w��K��*5}Vm����3�t �"K_�ƛ숲��Hp�y\'��q^ �"�ɣ��h��y������ih�.0�dL�ωL����6ުB��oH8�!���I3R�Ë�:yI.u���:�o�m�	�I��I�/~\[����)S����3� �ڤ�a�5z���gh_uRģB|�v7�V-���L�1�����N��Ry'$��]���w���ӈ���Q��Y��R�Ac�~���D����*囀����Cq�;b�(W!pT�WZ�(i�����IH�V���B�X#C�fVRו��^VPJ<�����:�F�]\Ȕo�2J��B,�X����JuXP8�_����7��Sv��Yv�� !0�Vj��H�͹��|M��W��3����3}����h��( �PH�!c�uhe�����ZZ���� ���Q�&�ڏo��S��FXH�� 6�鍁�'�q�������~�5kC/ڂ�
�>6�Ӏ��J�ܲ͞�Ĺ���y���c��2!��>?�c���ϖ(0�d��JƯO�C�;��Cё��/��n.�aKCp	C�8�]�k
����0�Re��?;���9�Uז�O��C�������?؄��'����O�-�/�g�7Yx�-��c�	��'��?�7h��b�H�?�����_P�ƗC=2��1��$���=@���M>e
![zt�{��_���0BjOyu`F93��(_,po0� ��Ս�E����5#��]��g$�7=�9�i�ag��ݱ�$�(}�x�H�cϴ[�-��uW?D�2_'
�6�b�\�яI����%3%5¿Ƅ؂�j�fk.(�J(
u6=G��<p<:CV=Y�������02�^�XM���$�rÖl^ÿ�;�̐5��b�ŉWF/*3����
��/b�q�K^��E�=��k@C�lo�Wc���?I���w����|���U2������p|06�2^1�"<�5�a��2��M$+eH.�Km��� Պ�^�z�Kck)s\�۫f{{���������A5"��٫�R�m�U��$�یz�j=�������3T,xk��'˩��/V�Z�&P? �y:������7?I�is���:r�Pγ�o����H0W�=݃��B.���������"�-�֦t:m�]yp�<W��%r� �u@t|D�:c�g ^ �@A��б�J�L	I��~2���Zla���z�ם�G+*ެx(`�l=��<O�����R�#�>/k\�a�V�u�y���ͣ@w?�ݞ3i�*�l�6��]��y7�*�ͩ��;0w�o�ܫ�����89$���j/YފC��`ĭ����ƀ�'G�~�|q Z&q����<��R��.�P��(���yT��ۼX�J�Ig1hE��b%O0j�Vk��CN�<x͈`Y�����
U�WC����stR����ziA�� ���璀{���D��lt܄oP��R+�u�"�c,(1.PV�r}#�
,?�M�o����y���QW� ����cPkD�
g�y[Jk`�W�j%<u�Թ�.�Sٳ��ɬ�*��]�1�:�,���(B�����2������"���=�����
%���%8��+�C����	u|��S} &y�d��G.�������G�[6
��#�@=��9f�do_D���3��1K� \dXAh���-m9,��=@�Զ�+A��$������N�ʔ��[�i�#�v@\��W�cה�
��h�)*���,i���UT�'h(�=>cIB
��o�XYr4�;�'�!��:2%,+�w��뛊��q������o`.�j��d!35��~��Q�r̶��r��^u�:��=���R]���Ċ�+�_#(~���%��#�n�����گ��i�,t�����(]���m���C���O�9���0zq�d��Ig�_qׯk�c��z�:�^?@����r�i j����Q�� �&���N�9(��fn�9���%��XW9�g�\)(om�K�a_g�\wT�*Z�8��͘\b5�`{%N��F�kG�i�uv�[��B�>3s������P@���W(�ϴ�p��(����0)qp�K�4nQǦ�V��s���%=�����_c34=�T.`c�xؿ��Q�8���QP�޵i�ٴ~yx4��.z[�C����,�#Q|���t�����N�1Xi1�\����#�)���QQ�p}�;I,anb4�ج;ݥxD��z�@:�����:Vˣh1����e�kVS�{g޷4cm��*N�{L��!/w�0a�Y<6�m{cc����X:��Kd�{�(��1%+�[����?#=|Q�%�8�CI9J�نiwPٖ��D=�s�?���"��^m��0"�g*�0He�(� l� ,��?��=�}\�_2it��Q�8A���$���N��� '��}�3^xC��ݺȇ��{�W��L����<En� �Z�ͪ��l&�q�{ԫ8�R1�LM�{}�ҕV.���N��?��qڱ3jhk�y�J��������?�d$:!�{��1h
Ś}��G�&|g���H�t�{7e޷<��w��(������AފD�l��A?��[&���M��e8P`� �F���?��][�y<�M�D8)�(�b�R1�Ra�%�-�):����J����w�eܶ���t)������*�Z���=�`=��e@�|����Ill��q�aE�
���lL�F�{��/�+�K� gE�ZHJ�J#��l~2�!�/���W#�:vu)��ꬖ�M��i�,�> �R�B/P�Ņ�Th]e��e��C�b%n��ݬ,��� -��q�!����#�q�7Q�F����X��Z.�:$Y�SO{�`{Cu��j�=b�q��5����m�I��V��щ�B;w�> h��#��BJW#gi�)�8Ck4^��}
ɵ �X7���5[���OD�=�!Ҹ�9�o��Ny2�pP�~zf?��^�����>ru'+�^��6��V@f7��[K��K��}��E$���54]תR�(��wM1v\�4�0��he售P���Υ��o|iB�al�`�J���� yF_w���'�ԡj�i�&��e
o�:���N�� �.~IϬL�m#������\�B���x���m8M7���ۓ����c�?���v��i�+�K��v�<��A���� ��$��OY�z;2u��U�s���465��;��Pŋk�-�W~H����"�!C�©���0/���@�����|�s����x� �Z�P�?�s|i꬐TD�[6�#�^x��r���,��Wh엵�֬���$����r]xN��,�<�>�&�xw�}�¹g`�2��^�_�B�߬Ƀ��2�V��o���Wˑ�&׺�gh�@&�kuW�VΪ�T̎���w�
�[��_����H�Kj�h?�I�:s-��~/���2�:څi���J^�O��G���$3,c[6�x&�ctj�Q�ex�����z*�Fn�.\�rGo���1ˏ'
���ܝʔ�<x�7���_S��Z��=�SC~`�8�rɊ�!��Ũ:+�UҜQ�,�����������%�3N1��!�{f���lfx٘Tx��3���J4�?����r����m|�wnP��C\�b�F8ǧ�?���!ߺ�i����hGK۱wd���F��X�C�7�M+l��MX��\w�MV���w���Rͧ:�̕4�#��;���i_�w$r�2������c��A�38l���ծ�NԈ�9yd�c��j��ct1��%�����Lq���i2[+ѽ��qtn���we�a�$V��,T#8�CʎA!"@��S��'kE|�l#2G�H���D�x� v�3���~*�3#�B
B];���djc#&�Ȇ��67��*M���R9���k�Tn�Ht��2�t~��E���(�2S��z�����<ZD�60ɔ�h����J����"z��8H���fXv|�Lr3�K��Gy����>/E[g��e�}
b����Xۏ�P\�M�D��S�͡
s�p��S�(��c� K��Q7.�T������!k7��|=�I��j>��uAadax�40nmI�C��a;m�Y���I���r���B���SGj��s�N ��:I��Z�$�Յ�TE�H��m��
�����^�F&�s��!��o��N^]!ys�զ[Ð�[J�لI��5�;|�y
z%��u$�;F:ͱ3�>y��VE������W�H��H���,Q&����@.;���CH|��ʕ��6�@or�}DR��L�	��?�B�[��N-�ln��\b��ԣ�ah;Pɫ�g������*��t�Dp�b�L,Ge��p�sx;5\*��ȗH��2>�a��Z#E�d�۸Q3.�v��W�G[sʐ]��y�G���C��@����;����)K�?����g� &f>���Է��'CP�����'����	�}E�'h�.A���MaP�G$�ARt��p��yO�j���𫪣kr`��g�Z.?�p�v�i���>M�ɸ�8Ac/b�'��ҭd�\xDW�p{�MU�RpT� �=�4,"˂����Ŷ���^z�&G�i )��F^ݓ���\Q�Ѿ�X��}(�c��S@�q�h�^ꋐ>S�
�g'z]6�����{4��U_k��'OZ�Ki���[G���
}�31Gv���l�,#�F���C4�������3Nx����IZ�e�X�~���S��B��jEY>"0hZ"������R�O���k�����rd��kd6��sGa�=�gh;��b����
�Md(�S=��̦�HDm&Y��b�4���7�8�l�����E�,RL�"��g�*#�~���$�,[z�k��H�gJ���I��*��,����P8���2�H��:��r-׍�J>D���ơ�N0Ne�Y�12\��`��<�2��\��
H}?�y-��O���+�wǀ��e)���/��m;]脥ֿ�ܬ�+|���N)X��:�=�4˥º��+f�#��L��bs�n�|�#����.Sр������z���g�H���w�N�y=JO�xeX��A�֏N?�>2#���?LW,��~���e�
r���&L��B�ʛhs�x4���g����3Ҷ�a���i�H��Ҁ^}J��.�%�s�����042��,�",H�jit��m�P�n2E���_~��~Ӻ���)K��Lsa��Y4qb�$�In2eW1��
�������Z/��X&�A�ٮ��Y�v���ɳܦᢎt0�."*A8��"���&�B�r*	~��S ��v�z�`'��~)?R���(ƀP[���O �9Hƺ���SI�~�#�w��i��Qq}�c��8\��\��_`fȾHB��y8��_��E�^8Q^Z��#��>����l$�%ǓKZ`�=N���x��oM�DK�W���KK��	�5����3��|�Wv���ޯ���KD�(ހ�6��t:r�����4����3������2�e�
�3e!ћ��u���$�^dF�3�	��w���`q�lJ:?�W6����v:k8�}����F<�Ȑ�����D5Fr�CF8� ��?jk�厢���.2���)���]+���5J�i�[;�ڮX�uv)�hW�-k��z?{f!�^��ܷP�+ N�hs,R­�?���o~��ݩ];�7�>,����4��B�W�Ab���m�$Jʲ��{ɓ_������=.t� h�:AZ������sI���Z;s��z��I�(����_�Z����L���DD:��?�D ?�ȗŶ�#�/I�2���,\?KC�"}�|��,������/>dIN�Q��vl�c�G~��Z_�3�E`�\�p��DY��Շ�Q572�_��I��w�'����A��ث�&b��ؾ!�f�p
3Yi9K萜`}{��u��B8&�����y����R���n�XƼG߉�T���<�0���l��<�~��v{f�G[�	#�.���I�٠�_����w|�trt�
i��c�ȳ��#����	���<=�j�Ȳ��ψ�Bj����NA>��B� (��M�$Sbu"ob�l���b�YRIk>�Г�����w�ܾC�
�u��"&��e*�Ɇ���r�p�$T����rJ��ܺ�D��=X��*�G���/�LDR?��s|�w�+9k}���/�C����;����V����)%� �b�m����U[�?]�꫹[��v�j���Wz��*/_HB�}\0��zz/]3�@�0&%�;���;�e�<j@�fV�h�c�O�`��?�q.����ih[��o"�ۺ
�����pT���l2Q��WY��;U�-ҟ��3�$xQ{�JF�v�O�D9�qyPW\��>Hvǯ����xM����zP�x��HT�OF#(7�&��-�k%�x�	 ���>h�y�F����;��U�b�6���������F��
AE_<���G��-�g��{�!���I2�{�2����5�Xq/5�f�V���H�[iB����:��1�����oH=��?�����#�w�QL�#o����Cyd���y��d�W���>�U�-ʸ��;��Z��=�=޾c���W��翋/��޳�By}��P<�%�?h���ǭ$Li���Q��ʵ��$F7�O��}5�j�����Tҽ�/���i�,T�Г����'��A�7�;u�9黵x���JpW����=�H�hdo��2j#�/�-������e9r�6Y����Z���h�ҬN��B�C�4Th��g�� OA�J�E�]_ւz������)M��4��Rc{LV�Fb��Zl�C�?��X=W��%�����R�p������Զ5���5���2��.�}<�
���+]��c�i���j������W�9�Mǣ�Y�5n-1Ȅ���m&h{�c��S%:�}/�q�܈\�q���Q�+� �v���߼ۖ�]��uD�[u"�y��(��U{�˙�/�I	�ݳ�h�/��zǶ3s�3¢��m�f$��(S��e��i�	���"?�m�"�U��KhT��R��!���l1?2Z[�sl� �B�e�x���1���t�j�N�Йc�����o8M#Y/N�����O=d'��T�%����
���8��)��%8�O�.��E+;^j�w�cU�:�JE��;��5U2%)�0B���AD2+�Pݰh����	���ܬ3*4�OJN�j� �{�L�u��xTn��[��h�t!��2/��y����eo�-& �5�!���i��.����rB�D�)f��W�ě0]X�j��q�W�Z�.�jBQ��We2JDb�K��*��ɜe&A�U�����P�g�Mąrw����pxa�����D������UU��.��g�����m*ҥq�9� �+#�����l���ޡ��x^з�Ś�}c�AU�u��^���մ�S������Xn��/~`k��ܿ�{F^ΐ*oNo-�����i ��A$<�f��Z7�֝��$�8~K�a N<Y�Ɠ���sp�� ��,�TDp�K���	Q�X��B�ib�]���uC��E$��)�� �@�^���
V���ǜd�7�2{����Ju�b�����X���lg�2Cw�fA�>"\�kLk͕Y��u3KN�7%�a�s�8TՎviVo&z rs��4�U�_���l���\�����[��\F�D痔�`�
G
�����-r�H6OS�0�:��P�qg��@�;����8������b7��;���N���Aٖ}�56o�aǢ�̤O��&Lu�5N��A�\�~Y��5��*��sO�'8��m.;RT���"�I<J�up���`�,>�
�X����)�ϊ0�Ts=�5e��C��X�#[CV�����WSk�˲���e��fv�	P���h#
��UuD`�6����J��$� �������jO�����Ʀ7��I~�c)8@)�,:k�ׂ:bɱ�ڱ݋A���E�������lj�a�U��b�g�5�޲{��,zM�9<k4ͱ���oҨs�@��G�R�!�u_����0��ް��N�Z�Z�~"��ű�6�b ��!]�pi
k�4����	j��}UdzÐ���FO8�د��\_�ʴBOf�A6\�8�IՔg|T[��D�?��N�xQ6[�]u��q��gݐ�������2�	�������-��.{���>G��'�)���	�	�{�����5:Kd�7G���MR� ߟ���X����i����P����l΋�/o����n/9��罡_̣��H'�ѩ
�G~v$5�՗V�R��a�wʿ.�}�mm�G�d����Pc�ۢ��C��͛����`l�lk5`����~�\�ao����7K��^�>P��Ĕ�o;��ɚ�5 �WN��]C��]Ͳ2L�v��"Y��A:Whs98%�M��'�3,����ڱ�yAb���ΠqÐ�Isر�F��e��H\���id�aµPx������<���,گ�qh*0~�CoG�S�%K��y.%p�;�R����:3ڴ҉�'��lځ���*މb�ٜp��ŏ
�̶���x.)�f�G1�[��ﵺ٣$��U��m*��H�镒�\�p�K̐�H]��t���'�á!��E��u Ki��B�#!���
�J��� Y�z���X�F@�I�����.$2�Q�Q^���(u��ۈ!�<'<��ŕ2Ks:M����R��-���r��i@���7�0g��j��6�/U�54�٬򁵾-[�!P6ꋌ��8l�
�Ƈ�[^w ��f� �]��'d�8��v���@��i9�������̏ $�� ��_,d�xa_s�w.3ij3���!g�r3�H�_���m5�����
s
YG_U+�:3��7�Е��� �MN>ݔUg���������c�����	g��1P�l�}������V�a�vi�f���B��][]5�U��dI�m��Yt����^�a8i[���s���Npu~}� ]���J��؅&ҿl�'ܣu�ؓYRl)f�
1��N���nzL�Nb���`��!�E`����6/h�`V8ǗQ*����OqIꞠw�EL����<9����,��)H뻷�9�s-J���2��v����R���ɒ|b+W��^K����G��1v�ȋ�_�f�yK��Os�>7�����%��IT�	�{�P���_y��>��w�X��9��<G����u��^���t:(�6�; �Ջe�yZ�HRc,ڋ'�X�E�+�	ZY{��A&0��x9��Q;�l�ƶ�?�F$��'T�*WUs�_�*!��Y��Fr��FT���X�ֶ�r~�������O�v���O���옺</��Z�1�H�Z7�ã�y�L. ���m�8��WO�����4�NQDN!D�wW���G`Ui:��jK\�|F�1u�s���g��r��473E"$��B�_z 1�>�w��,t���@G���+��:��^t��qX�����|ɮ��*o�̶��{���B�g���Vo���S���w"�·��厅�U���ޓ%W	ԛŕb�Q홱9i^ ����0$�'+y��[�P�
���GY��y�T����=��0h/���q�*]�a���]pJ�Z�/�x��l��?�g/(|�$6��`�X��!ĥC��6���W�r*�����M�`�^P��4`�ni���)O��!���Lf�Q 4�?�7�_]x4�׿�y���|A4��m�&�T���4$:�6m)ѱT���<��	�!ҪrNy(��s�4J�Qgo=�5���^fgQ�,�a+k�����!��.+Z�EJa�A�����>˹x�bW���%�Hz��g�VL�Y������ƓŜ��,�hc&[��S�V67��x�XeT��@�%��¥*d����ܷ������+�����dږ��agL{�W�k*kH��K@I.a~i�jnjO	ᆞó!2�FY�̀P�Y.{���q�)B|����M��l }�S���)���`�z��غA�O>� N$��m��#�5���8�q����=O�
���d����
�Θ��P��Ը�m�S�{:�d�����ߩ���X�u��Z�֫J��^o���m�u)��E�Lh*<	���Zɮ�qK���PSW/?�Ħ�f��iG�Wx�� �#v e}����zǃN�B=:�L��L<k�f\��@�&Ʒ\`�mkqf�܉A9� ��B���ϺX���[�l7+ֆ˾�:�[����.��c��k�`X�rtw�¸�D���<�-ׁRc�V�8�
�͚_yi3E��3�մ�yQ��_�>��U�xN���_���7��.V��5�ޒ��M:�1{;��K�M�P�Nr	HfN��.�gٓT��h�`��0��ʆ��nc[^fZ�&*[���a#V�I�<���Dv�Cl����ѭ9��=���*�WK�X�
=�{�G9�A�U��K�*��Bה<>����w��k����i}}�PR�YX*���@ip����Q�T^��� �5���E���i�b��O;��ֿ&\)�x���'ɔ��/t.z�j�}��ݶ�(l��l9���ѐ�V_وl�j#�Y}ETM�XQ��ls?��I쭼���U��7�_��Bh�xm݄y�4z�R���˫{�ќ>��!��t�Jo^�_��#��d{������T��e+�s�Ӿ���Þ&=���X��3�u	m!����𭚰ų-z�+�F$տ�\�U�v���۞=F@1D-	��2naa���B��g�?��J��S�k�I_*��ؾ��M|�g�Ԙ�C��̼� )$�I\V�b�PI_2Pc��;ԯ%�����Z�i".@J�+�N�<8��`�e�
�!ׁ��M|y[�$��n=O���h��+������k�JO�-���EUb��Yv��}X�p{��|{�1��~X�Mi�^Z�C�c����f�ZצӺ\�4�J��4��+�A�0	�L�N:��Dݳm� �E����.e�Fq��S.��t��h�W���D��~G�F9�V��MA� P�ғ4~� QTB3�B>v#-x�iW?4B9`�kct{�؝��A­-���V��T��;�cff̲3`V���L��UО���٘��7���H,�Z�T���L����M���V|�rz3���1b��ӑ�_��vр�]m�`�%F'cw�K�}�ӗ�s�:[�SaL1���#*=Sb(xR��?�e�[`V���^�p�
��.9�8��U���Tt/f���f_/N��1����Iߖ��Z 8�5��$�O��
�^�tc�7�8(�1�d�{��<Vb��e?Ǌ�{�$V>����q[�	cK8�%�����g���6@�@!e�д�������¡*����B>��z�X�+1O,�He ��>�~�?���{��Mp�"WH��m?��xu��M�?&
c��Hf���;�G^�pU����{h�ڎ���Y���E�VLM�Z|��_��-���v��\?W"Ƒtp��J��0���Հqq���H4
��h&�7��ê�%nx��G�/��1��-�V�s�>ټ��^���?��. �}�}26ck�s� �ihB�L����X�nfEqd�7'3T�_y �7P1V��S�%��%%o���N4��J�;���-���1�KN������"��RS�m׮ة>�4�L�c�0��^��>+�*�p�cH`5?^��Ҳ�Re2^�A9����W���ckڿ �{ ����dIrT�D��@�2���?�(���7DN��֗�w�nKѽ���1�|�H�י�E���j�oW�0
��c[y΍����rʔ�>j��M�|i^J�s]>��>.ygP���P�y�8�O��K��K,X_��]ov���+�R���y�����Y.uK+.O�Nr��kɆfRL�j	;����ߜ��Q#evg@J���+cV[��#ʴ��+3fW�J�0�|m�k�� �}I�����e����U��yC��z*I�<��$��M�ϘnƠA��=U��w����H�xi[�F ](:U��E	{�'���H��K#�I���]���6^�����
Fɚ�7��%%@�P��-�ܻ�I�9�^�X�w�ү�D�����1}D<� 27�I�W��4�(��w)!�H��j�anŹ_q�Ad��s�ٗ7�t�Ȥ���)h-	�"�L��u��͂0�Y�����^�N�'.56�P�k�fuA����m��f�����ND�AkҘ�����5��z���V)���o���G�#� ��Ff˯XF?~A�M1@��<a�-�:+��E@��h�س�2��>��`�	U�w{��X3����A�]��x@���5�Y�B��2F��6��-���لY�&c:7.�^����o��]��@��qV�_��n#|o��ݶ��[�M��_P�C��%ɨՃu����U@f���dJ�b���gc��X�P9�n^��G�ÏcD���R��A����o�p݃��T������J����}�G��:������:\���m�<[7�����ۡ�@��4�Xm#��<�W��ֶ���@��LtZ}�E\9��P=x�W��\�=�r����A�k�)g��~��OZWR�|�Y`�����]��o��I$M�)+���zuj.UH��,:�N�h��X�M�d5X0�Ժ�����\J�@u����;R��;}g�����"W�a�VG#1C����3�jq�����?"�$v��Ej�W�d���$<���Yr�Q�<͉�=�Q��%�]<NE��c2Ëo	(� �ЭP�cMέy4�����Ե��qIwk~�Z�w����:�}X�ʍ�Q"������	M��G�G�ť����~���-�e�9�v������&��Ż��������X>%���!ZP<'\r=8a%*.u�V�W��tb���|��ezx�Q?.n'=x�F��J�4 q�Ŭ1~�}Ŷ�1�A�I�%O��z*�w^�k������ϐ �������C!]��E/�aF��J��N�~�9R�����gy#]@��z�����p�i��@i`�hpB4p��\�q��T��D�?¬�w�XN��/�� �{�J���es�}��X�"?���%0'I�^3K��~iĠ�ņ����������E8M
��N����]�NC�
���-��E�>���r��8����O���g�GS�Ǉ�ǪL=4ހ<�\K��H�x^"��#>��k�q���0�_7�'&�ɸ�⓾WS�6*��X�Q�>�{,��O�_h�"�9l���;��R�PگEp�E)�+��5�|(0��@��C��ɿ-����������eՀKd�;��ia����~����ĪK��I,�=��/8d���Mµ^ĨR e��;t�)1�~�-�� ���"KRR�1˂l���K���^�n��$���?�߫��q�C�W�]}%`�X�����(��!,a��/��˟�ޠ��p��1'�i���A��P�:~�a�%��m��2?S���������&�BaD�Yr�<7�Y��e�������d�I3�����E`�_����QMf����ܬ.��0��x-�Cg�GQC��3�I��S�(�̬���V�a����(��"��?��)R^w��Ï���2L���[{o��'z����h¾29�����_y���ߏ��ϯ��Պ5��5�Xv�-�Ǻt�j6��N��h�X5��ݕj2��K��;OlW�%N�WǓd4�_��DCt���l�ӰGyS�K�mF��Z}:Y��o�R� ����f>���t�����.��
r48U{�o?ź���:�41f>9�1&�G�'z�ڷ�T#����] ;��O�!8ztvʽ�?�e)�"���=M������	x�T�SZu�ј��\rܬ��ÉS��(�sA�J��J#�8�������K�����Ԅg!*g��CT���_zD�^����Q{T؂��ܕY������"q��++��-�w��� ��a��{�����bkldS�;��٭!o���\�3�+~4��'Mx5M�����^�O��ؙ �$w5i��%�-FL�����DEs�h�9��l�ֻ0��#L�a�pUR�8�K���hTB�=<�X?�5�b������-G�����y�}�~�ć!G��9�Sk>M汎,�9~7&mk-y@�6"�x�zVjL�w�F���(A~�Yv{�Ҿ�b�@��g�w�ι�q3���Za�,��k��y=$�@�x�Q�Ec�;y�=KKgG��~!<)�������6��s>���ە��U)!!�I7B�IN�aQt�vÑ-�s{
W}���G����S� �a��J������k�I��1_�WnP��-ʃ�����Z�B,�p�7&	G��lȲ9�x=Y��@,��"+ΐ4~t��1NN��p�WP�?d	㯜w,����WT{p�&w�f��x��V��7���z���WrL+�L�(Hé2�i�����n5��E��ƚ��S"{@��� ��G�;d`�Y,+:��/'�����C��ؤ6w(|�.L�S�����A(�C���Qb���~�Wgh,�r\��.�_t�^X2��9IP����_��|����K(lXu�*�@��*��q����.�2$/ߠJ�
���y���ٖ98'�T���n<�VM' �q=Y�h?]fF�&�6�y���(��8���:1�Mkc��!�f��a�~י:-�y�`ޠ������p�%���7]uɣ��ةu���~gY��L��&�zz�QO>�������=}��q<���K�.��s��$�L�f��\����'_�]��DA�IW�B/B���K�O�I��������������T�%v��y2�Uh�=$�+�a�`+�Ln,C�7f��Q?�����wc���z<9�n�V��x=$��F��&]� gJy(�;^��Q�w�1&%�}h�Y[IcYz�ީoj���FR��\$>!����u���^��c7(k͑`@h��&<(�gD~H�w�;E���`���>��[6��1* �q{���W����E=*A�엓�Hސs��cȣO�1(U�0G���d���%�+2��i�5cU��>�*�7/79k�.'�sE[�v��戴���a�5b�;���α>o0\�&���8vу����V�������IȄ>��Ր�e&�6��-u���Q�Z��U,��8qAݓ/���+ýt�v�#iT����}~����8"�Z�}�1-��fG������R��
�ȱx1��6�
���N�ÿ��x~�I@I�ڋ�9�f��XUm�-.����ϛ���)����xg[&�\Aϴ]+�@�."�'�f�Mrj�����nPǚ��{v�?;���1�?��Xe��,�%X��9�#$cs�U���3�ԭ����f�e�>��}�TZ~-� �����F5���������q�J:٠ʸR������TFG���~��d�n��4�Ú�Aq�f��t#�v��L�������th�B���j�Ŋ~�R�������RtC�@j=x��y�G@�v�) ��ִAI�"c��a�'`W��
�(Vv<�� ���/AǮ�i�	H�I�nW�#�l])G<�%z�~�|�7A�lX���}��.��~Q��޹3r����4}���6���2;Q���';^8�,�B���?�w[B��:���[���z��퓋�q�)��y�-7/����i{� �����䃬u�b�I�l�ԯr����5�8�����[)��yj���{Mג'��q�k=�U�wc�5�i�=�Ģ�gZ�����iMb�M�uL�=���ￛC�f��G��Fs��~����~�,ä(���2-�pD��*��=��p��3�Ԗ}@Q�]��E���rǳAl�67�a�:)�C����Q�o����[���L��k���ܰ���_� ��sG#�[��$L� ����T<�)������\��1B��2E"��_��X5�~*����P�:�g�2ǹ?����^�D>�El�5s�a�ԍId)7Rd��r/x�m�g���}���r�lP�1���݁^a����~�9��99�Δ�5@���H�oMO��Q�`ങ����_B%@���U��^�є�8A8�w��`SbY�TA7Q���#�|5)��g��%�����W��9�ʢ�[H#�DI6'��Ԡ?d��������F���q���%F�=��!�r�	[�Ev�/��o�!��5\&��������C�V����'�?Y庻\<��H�'�O��� �,$��f7�2�H7)��s�;�MV�N�e/ꦝ|��8���O����	P�2M}�Vc�{ ����XP�L����S[v�FU�T�����~��7�Bx���Z�y�vև��G4�+L6�с�E��r3XiX�#.g�< �IߨK;V/�� ͪ���-Ӵ�5�w4��c���dM�Y�X@�߂D�h*k%��q����}R�W����d�VW�-gXHQ#_���~�"��fKZ(��.��̯���@:"@�b��e��ؿ	�i�
Q^�X�G�GS1*�VԇWq�;�!9�Q������z���z��%���w��Ns�N�D�%7�Ӵ�)�eW�y#4��Z�p���	P�ն�F�Vzr�J���*̡���om��R�N��e�;�:u^T�y���EHj���zŗKjPd��Osl�t�?����r���n|�O���@��_��I҉"�g�]��^����E�>Gt�T������h�J���"�&��*�-vN�P���\<�% M)�,i���."D@aĴ�C���ꭓ������$H��b�h��S��w�J��%�ڀ���V��gW'$�٦ԏ��R���{ksai_<�����n���w���+����:���#�ʄl�a�F
����dػ��Z�KH��K���|�:��a0����0��lQ�����]>Dڿ����+Y�l�bL%q�2�un�(y����ư��ޭ��H|ZM���|B�N�3{�*h�}���,��]_f˒#�=}����$ �/?L��{#��G��!��T��?P��^�8����~O�}��o���v�Q��-]ܝ�S�SBWe�O\j�_ebR�g<%�{�|œ`�dj�8��[P���߻-�]���B�5��nܙ���1����B7��ϡA�Xǎ�
>��R%;pelq`�9�k=p�B�ٲc��*_�l<�b�U����W=H<0��*��Q�B8���'Su�a�������YBLD�I!��	�A�����u�mQ���K�^8�7��g0D���"t���e�����\G�^�|�͏O�A�Ąt�Pm[������NHJ	�Dm���
��m ���\��_o]^�a�H�t������
?��|�'�VW�_~�*Uw�b|>	27���1�"lmDm����hkj٧�^�4�-p;�3�@N�`ܕ��� �>�sڵw]���d ���s_�ڒP�
]��. ���6��71ƞ�Q��J�;y��O���xߐ�������w��J6p�(�����A��9�r�Z�g��U�i|ٛ�'ز��br� }���'��h�C�ź2��Q&Mh2yZe�R��aZ�8�4
����������:���ƛU�h)~��_<�
%����	+t��	*S���.~v���8Ew ����pۥZY	�(�ݤJS�`d��N�d%��
2�	i�gd<�M�Q��N5�*w�4XDb?L���'�#;s���������2�{����q���7��x#���pH3HT�ܱ,2���x�Cn���<���B�=�W$���5� �ހ撬˨�	��<@��!� e� i�w�6�p/��F�);�5�(,x%�X�j��S�!E�~oE�S?�hy���W��P��P�u�T�1]L� h@��ЈR������V	lsѐ���y���m���|��8��T�noꄲM�d�m�c ���]V�QXɫi�@�ø% ���K�+�S�s.�/�"�c'o���1$PKĆ[��3��ЀAbb�|��+���Z�<ߓH��Wlt���f|���SG�B~�H�A-,���QI �W�V;!B�m�ɢxI��r�O(�����S�%Uº0b�>XՉ��ڢ�X��w�Թ�_�����7dW�ѽ&vjX�/�v�^�Vqկd-X�L��3�^���@9·�Ig1{���:��0uw�3��}�l"�K׺|d���!��J/z��+��RVl�"���w��i6�x7?B����g�Jc����G��6�}���h8.�5V�.���3G�ŀ�"T�@�q��x�V-���1�:�D|�������'��m7bf�b��/x�o�Q1 ����[f��KwM(�I.[��&���2�[�}�����xeα�m�s��R�ej��Q��@��_Jg�o~��س.�Z7����q�_�D�E2>�)�RB~Y���X���	�����P�
ϡK5Y4�X��\���&ҩM��߻�2�2lܭ��<� m~�NS��S�rkeR��w:��*`����K�j�0�+l5֩�3ֻ�=�������m+��~ӤjI.~��N�p;)���S�3���"���B����e"����qm�~�N��M^����9ߓ�=��w,X�6S�S�L�^"F�/y�8����-�_U��M^�4��݁S�b:���6<��֝�U�2Z�q��.�
y؅�Ŏy�!�nW��_h'Z�k���}��������������3z9�o5S�>ǧ�9��'�m�r��1�ڴ������L{BW��fN)� �B�� �����ċ��ю[Ā?Mѹ�E�Y�D��������m��x�q�:�����f7����
�ǢRg*2n�H����"-��v����Kp��s����$|�ɒ��3�>��^S�N���2��?�p=]z�q^[��A���&ƿa^p�2I�������r�G�x��8X R�b�A}��ϲp�\/���=e��F4y
�� a�����h��c��DU��~�m˃-n�,y7J� �]m؈\��1Q���~��6&P ��A��A?�������_/͠9L�v'�kn!�gq+��,�IQGC�l��,�c1���N0$ ����J�`�y_�e�}�s�	��2J7��%�#�|��hΎ>��G�b��*�j�	��yr�s��ٲ�|��n`��J��3�������f����ҋ���(#�;����ύ�-Ql��!��?���ʍkC���D^B��v��x�%����5����9-I���<<8W��ND�h.1n�כ���Xd>��yuB�*mBOm~�{o=������G��P�GR�Z/��W?Bdф�%Z��N����!=[�:��lm��GִI{Ͻ��4�-��-3�P��Ii��%$�xB4 .���,�K�� s���$e>Vr?���HW���c�a�q).J��q'���,���^(؝�+	-)�w��NЯn�t�Ɩ�Q�U�ǯ=e��өGAfNDG���z�l�S� 8B~A+5���!S���}s*�����a#~(R�&
��Y� �잏��{�U�,�x
(���%?̈�/@��T�����u����ʍa���B�^�����Zʻ�㦍��/��%}��-"X�:�I�� ��ҝ��6I�����V�J!$�(,P��b�a�pԵE��K���w-����t22�ק���yܖ�n����s���Q�t��P=T>�h䁑��W[���f��}C~���JI�2S5��C�Dk����/�օxK��P]-�j0�7���w��
�AM�-D@��zt�=B�H֛W1z<��%'�ǲM+	�!\�v���	�7��
߷�c�"�?D����LnA�n����&&�|2\^��z�$M���~l���/ͧ��v����O_=^��h�3�:;酚�b�Y��#��,����j�����r��^�l�
��`\x��t�!�mr3�N�*�������/ܵ �}$����ö�cE~�v�զCxC�s������K��uBO3f�ҵϢy�k�q�QE'nO��@�v��"ԙ>z�yI�Q�<��� �M�9�AH3H�M����"#|��r��{�����*��g�d� �bER��'��:���-~�T�^�>i������5G�%k�r�C�B"��r�g�?p(�9�u���{�e�;���t��A�SF��:�1y`���ZM4��v�X"Տ֥ٜL�t��c!���2թ�͢�Ơ���ﾋ���FB�0ȒvET{����=�ے�z舳ռܯ%��F�/�
\&6�5\�A%/���-���.s���1.�C~��1�Q3M�w�����d����sl㥪�2.��iǬ�z1���ɧ	�zw	����SD����	��`'j�iߔ]�u�s6�pu<[�>��/?�^Zb7n��-9�P~���*	�?b�w���á6�Sz� ��J���N�:�G�{�+%��<�`'Il��e��_,�r���b
�T�m�?}��̪���]�.fN�vx��J</��/�x��*h�s�Jq���ޢ�ZCZ~|7�T� ��Y�RyR��ڔ� �L	��{N������ 9q/���\d��w.����p҅%S?$�sr2XWBf����
b�6F�6��*�V���>D�i;��M���p��Y}�����qm0g«���N��X�9��bg�Іo��N��
�c/�)������>����nY:��s��V�1Ԕ�B�{���=�>_�῅֠�7mn�A����iB⁗��`�NVg|�8�?;ڔ%y�!b>��g+�+;�?1�C��Q�4`�x�w�A��c	���|"��(ٿ���M	*[s���~c`>)�SY8����ϯ�t[�{|�s�.�Y@��HB#���U*��ٺN���,��0���C��P-��yYa<Mw�],_�cbR�����W��o��,���Tf:d/z�W�Sb��qPn�O,��7�w��d�����vc�YQx,����H6�d6]��h�?��h��W{o�ex�
��o���j��d��*��_��
���l��%{���x1M�'���@���q�q�CEw��p��l	�`���e�e�.W��ދ$�G��G�����N�k+��0�nq�R�`�SK�O�������Lf�]�O^��)����k�ӓ��"�� M�a||^Ջ���f}$�;L�2Sy����.U8��]��5nԌ�N�!h1�II 16p�u�G�X5��i�x�3E��!\Z�}[q#P���8����=��'E�,�h�s�![f�ӻ/�>�	��4�-T%����h�Z��zBW�zL�H�j�)����3�B�u��hvl��G�����yK$ر�\ZL3���Z(�R>�d�w���~�z:fò�$m�]�]#,�.z�9�B.�A�Ͽ�;頣��������$�v\*�W�َ읅��+0��bz��:�H�M5�k��]��6@��pcR� "fLZ(�t"{6��V�z���z,�N%��9�$��W:�n�P��,�A�\K�m//����'ek�����!Ȣ�H�Ft����������c�=�ެ�ɪ���p<��.�:i
~���H�#��Ǧ�����{����k!�l�M�(��;�XJ��yEd�ٶ�w�G�>G3��!X�W���Z�Oç9��`y�Uo=[�<~P[(�s%��4�*�9k�.]�������^c��ʔ���즬nVC -ܭZ�2�$��'	Ø�u�!���ޙJ:��~L�@J���TѮsc��l0�i�~�B�s'�~�5V�L�&T�f˖������׿�͙��={F�x�c"�S4M��à��ύz�6<�>Ӕ�sKL������_%��L5��x�b���)�����>A���%<u�V=����^Y�'� 1�Х#�D���X 
H �DA�"d5�Sa������>�Z���4-��H���w`7 ��Wmݏn��6�>p�}
��=C�����1�Jb�'t��r���0����,Q�K�w�4M�R{����h�]�VJ��|�~0�B\G%�(%��9+���|����9�4�7�t�dC��@a����6_�v������C������$#ic�:��/	�L��W��g))��Y�:L=�ǅ^7>iwz�h�@�R�\�&�{.de����2:��t�Pr�z+�eX�i�j�B��W�D�>qΝ?���}��`3X��
������D0w}��=��M�a�!�nϬ����i�#�u�b�K#9�x���2�8L�e�_:�aXY��T���R3�fS.5�m��ֲ�^�['��d	�\�M0��A[\�cx�9m![/�q��o4y.�o�	9��m�C�oqA��L��lO�W����B^1 ��0����l��=�09�p~��nKE�[�)��n�۝�?�MȘ���,0ȓ&C�(���5o��b��8��Y���V*�$�B)�����9�s�yg���Lh�V��0	�����"�W�ŢEƥk^��
]�2�J�VP�n��B�`;���#�Z�{8�r����tfl��y ��_��e�C��BJ���?�����YA8����v�o�<��i��R�B�I='D����}�o���k�.�&A������YT���nZ�?����o�#L�+�Q�~Ɗ������,L��^�rE%BhT#��`zJ�q+ߑ5�K�*]�=�/�s�H��V�4�eN�ň󶘟��θ_�Bl	�i[���c��ޜ�D)�N�r��U��p�sG+G6�ф����A���;쬟�GV�Q���c=�kᑆq����w�H"6�J���eZ�*�ZPQ+�����^�8�	j��-6<�q|��K{}�`����G�C'q����1Ĉr<}3Q��o��A����G���~VK�Ŀ���@�T��=$��ʎRR?����/./����w�Q4�jA��I����d�,.)�K�I�h��Jp��E���e?�Cx=߻��VV3RBz�՞�s��%5D����IE{Zڧ��k	����>�ű����^e)��,���h�Ȍ��z��/+�{��Wp��B�e�wx{�g�{V<��������=ͳ:����n+�)VZc�D%<�z#X�[/�o8�
�G�$��ļ�՞9�<�3+ت2ho�t䕼�}�1wjP�qFi�S�:/m���W�cC&t9~4����<����>�JA�.���W���,�+�%H������9~d���f)���?a��}�P�K���v.Y[�='
Kl1-؞��qQ��p5Ź�
	Or&�T�x��M�޼�|�� H�9-q��)�l�X�2�JfĘ��;�5��s�m���5���E�b�OC�w>��N.�l,0z��)u%�4vm,���d���ߴ.T�"��\���zVq#^!�6Ѩ(��_�O��E�4�',�_��AK�,c�
cY�i�t���#�FH]�eB��7��)�T6\�s,���S��]�9��Tx���Cg6����{dd%Zd�l��
$\�h�X��	�{$�j ��5<�ɟ*O/iXݧ��5�M*�֥��/���4Y���0�D�g�����jL=�eoEus��H6H���w�"������k�t�c Xqx�RQHZ�3�u��8����V�8OM��cmd�W$����?�{��-��B;�wr��!^'/�z��J�W�1��g�l_e�cֆgG�]�<j�`�t�ƨ��;��=.{i'9&y`��Ր��O\�"�2�Pŏ&���Dȅ�jFX�� �־���p��v2ۃ�!y��E���`�ʧk��������#́g��t�h�hqj3N�)��3���N���?�Z%*�pٻ>+O�V;���P ��ܩj�O��r�R�k�N(rZ��,�+2�F2Z`cߦJ}wh�k}f����uH���.�7Ż],�����w/z�,�v:Ңka{ ��1�P���zn��6]��t�1_�>��rj�	uW<�	8$�S[P�׎r�N�R�v�ψ����$Դ��-G�^=�J�eP��q�ٟ'�Z�=����N�I����niZVC��j2�WT����Iʷ�F@j25R�y���](�*���)<��c�7܅x���{k�7'�$Hs�Q�yrf
v}a���Ko8n�3�}� �oo�ap[�x]�ſ��{��v�S���	���>y���;іk�N	�y��;3�Y[Gc���S0��;�՚̃�P����W��s������]޶��J�lO���p*%��
�]�UfJ�!C�����>?�_���,E�-�hzɯ�Г')5�9�@|{]Jצ��[�fZ����y�zB�5O~JVe�>�MfE��ўd\� ���.�x�pWy϶�jP�B�탠11����a=�3��}
Jq+ޞ\�7���P���-.I@���,�
xN�1biA|�͵�_B9e�bc�"t(q,���w!fz8U�n���-{�ud�� ���t�#�Wo���'9�z�Aa�6����='�\�C���\�����Y~��`��l]ߌ*'sB����������yg�>� ���m�r�_���; 
GhB��+~!��y�����c����uq�}V5ԑF)��رw<Y]�8ˢ�లJ��ۋ�4�R�頢7h=�,����);ǆM�Au��?�93��=��^�N���9�a[�Y�s��=�A	�&���J`�*��ˀ}�c�(���䠱_�80k�R?�1t�y5s��D�P�S-��lAq�%=�d�����Q�|*R��L,S��|�W����>l�!�J���Ͽ0�h�Dv߲������[r�J>��s!��T�Bڶ��#�ޛ.��!�� c<Nk��d���_�
zki(.�C�@9����3�_SS������(���IM�T9��
��t����R��
�kR�?JF���%OR����W��b�]Vq	RD1�/�Xr� �{葾���/��1���x}�:�;�8���i�1�I����$q)�|00�=n��5�~��OE�O'P��_��m�;�V`iy9���c%�q���}�8B�dڽ0A�反˻ �`�ͼ����2��'ڑ.�V�{�b@)��jq�<�f%�ˌ�:�)���)����ghh���K���[�,F�y��}�\��dv��s�-Հ�3���ֈ�!��^�f�U�V�D�u��Za�e��n8
:��dIM]���l��ks�vG���)�d��u�U��d�� ~%�5_.�|��o�YbNo���0@2C��>�<�Q�t����ubo��=|~X�W�BV�O�80��q�b����Q|���%���P��"�e�YƟz��"(��#b����s�jn�l�TySM)O��zϙoS6U��Ҡ���U���>��N۟uEIdF*��o]X��� c����K�̇��|�R��ɰ򖐩�pJ�[n�Q��CV��7�|��4��a�dxNޕ�?�H��'�!�_
L���MP�0�.Ѓ��4�?���L�-P�1�঱D|4=��v�˥<u�	���7DV��P��K -gn��eL���ĹK`��W���̃�oi]}�Ӛ.��82�`�(�vM79-%�5О?��5Xjy�"��b'�a3`Ab����W\�� ������^�ߪ��kQy��`
��2�U�Tp���@��[���MR�Y}L1�݈��Y͠�
4�C-�_]����~ڽP@fh�A��ȥ���TD�>M9]rf
&8�m���O��N��� ��V����nm���N[O��n�O8Oє��(������G`J�~�j#�)�����&�	��<�?0Y':S݇'��(���t���˱�-6j��/ Ă?�r���@N�w�_�>���~Z�]a`<3v{tfM����+Hsi�j���}���<�ӽ��޼�ћ�qD%
�g�E��1�"�/2�=<3hԽ.�~��]S�Q9�
�`q���R�lq��*�w���E<^��C�Bc:y
���wi����d_�G'�}�N H� �K_ %�H�$	�C�Jl�C��5��7�-�2pMQ��vC��<8nw�%4$�F�`(0?(��*�.
�6�����D6��a��*��B_�Ny+�7��Բ&-�H���0��E1��@�
�z:V�B�)�ڙ�/�ue���p5]�x]��*,õ
��.��?쭆}'� ������:c<.�T -ͦuL�G,���VzcX�u���DEߧ�X��g��#���=9��l�ڝ�@DK�oCɢN�`.k�L��>��]k���EDf1/O�)�-H:4���?��Y���7|M�.AK����p��F�ʐ@k���T��!�Qv,n{:�kC7ժ��J&-�Dw �C��2e���b�	��&�֠`��<�� *5j��"áI�U�v��7L�q6�b��VG0�;����]�-9x����/)/�\l�s(�}+;�SB�<���h���*���QX]����L/i��d:�pWKQ�D��p��Z�)so��"��ڂ��Zg�)u��6�)Ap��N���<�������2�m��Q��9'��ڞ����`@����c�P�2u�`�hs�D�'z��:9��@&�����H�͆<�yo�	n�7�Z�����dK��8z���6�2��l�C6K�$mW�2�qN'P-QB����O���Φ �'�A6"�Q�Y�	0�6HH�>m2����|ܝ:٨F�[��Z42HBg���@+�o�m=��Uޱ�����ex0
R6�Qu5���̊����d'������3d�35`٤��'��[�Y�}��F���k�͑aC��U^���Z�' �'(��c�:Fn�����*DY���9��h"ZiK��u��FpZJ��m:�\	�
@mhqL���Ա6���d�ٟ;+�1Q	�p��u�:d&��hx�Y#��í�_�5'��s��,D�|j���r/:������#)���T�E$�ja<�f�����$B��P\a�qZ��"&����_�x=c��~,��M}0eO7j��zm��I]����S^�{�웁$jF3[]<����_�J���
C��u��n�N��ƨ��$�:���f$>��>1�~����=��0A*~�!���F��>j�c4�_������L�xO��ߥht�O�|�����~�Wڬ��חN0L��t�*.�zr�b�S�������/�?ut�)Hq���#x��?I�g���5��<�����F���yS��:!�:�I�����q��y��.S?;�� zj \��r��B�u2=�r?�^0ݙ�^$M\Ң�Ε������E����{���&bv�y�e�`�u�C�g�z�����[&�[�VEΙ����5��x �+���h��xbM��Զ����2V#�~�L�{+��F���WbK��Nd!��kGr��b�$���׳n�~�H�HI��f���Nc^<��C�� �T��u�����)�[�n�YY�jl�Ƹ9�P�։H�ܞ�#>�U�s, tu�?fF���݆7���봇��Wc�4\i�ˈ����k���%'h�=�$���iG�DËJ�3nW0<���Ws�a�RLb��,*M#���wt㊘��R��T�< ﶙ@Oh>և����Zr��t�+�d�����h�+p���A7k����Z�]�[�9���h���P���<���N��R|��Fx Q��q�|'� q��(y��yP�(�t@�Ӗ{�V;�����r�X-r����(##�E-��8��#kk��EV'�ՀHP��Һ�\���0ޮXP�so�=2���RW$��2i�{�s���]�����
�w���j:�=�mA���/�~���@q�T���2��w����nr���/�;�J��̖6k�c�48�C������l.�V`��`���<r������aU�(�����7�
���p�i�"%/�MJ�i��B�)� g��z?����澨{3�p=�o�|�_�5#��H/�x�	PX�^K%� G[�o� �#���^�|����8u�;����6�~����Db6���0�;��y��/)����몕�G��?g0MSu1���͡J�l�(:B&f }&��"�H���h����jG���^8�/X5W�zk�zC��EO�����V�eb/PĎ�a��\����k�=�6���;ʞ&���Q6Q�����|����&�K}���\����1��oP�(��b�6o�����`�������x$�K�"`��o�åW���#���|���4��Y���K��;sh�����ꢣ�(tk;���./���6�Ԑv�cy��t�R���
����|��v��G2�L���L6� |���l�R��4A<�NG�TFW��`	�Ħ}2��f�E!�Ʃ5É��{�3�?��6;�(+ÀuE�1%L��jFI��FQ�1ǐ6T��u�|�
0z{�����:�sp�-��돻�">�_�e�w����D��DiM%�j(f������.�<�{+w&��"�s��g� 2-���"���ʱKZ�%jol0����|Fv�����T��8�����o~��cB(�2�]��q8��a�?�.6���źo�)�^��1��2_+�h�i亸!�0�h����FK�����!�X�9��nH3��V�|Lt��Cq�V��+���}�)�J�7t�E��7��˃#�ðA@;���xs`u���O�7R�L��N��	㵞�~�āb��'�.	 Ɨ�V6e5�v���µF�f���3�K�}���������l�|s�,jmh1�W�k�zG
e�OK6\��� $e�'�#sS��i~-�YJ���C�����	�CE��ɾt����:�/��>Y�?kӑ��$�'��������T��vH��OH�z��&6LyG����W�ܙ4D7TV�Ib۲+���Y���1�}06��}������d�P��%�Tϒ���S����A$�d#���r�_�g�B��V�Z����>E��{�o�p�`--�e"Lj�ٷ��&Ӈ6uU�{���d�K"o���� ���A�{���������I�S$o���6�,Mк�\�9����.�NR*%{`���_�k7E�'J�nGJL����~�B��� o�Gۖ�Za�H}�3��
���=���x�dy��Kidꄆ �H�D��P!�C�= �T��z>�$��w����2��x�<R����K�g�A�[�3��>vbX��d�ݶΈ�+�8�<�d��e:�,�����mvڀ�
L��*8\�@d�5����P�O��@4fr�fp��2��w���C�_�s6��v���N��77�e��;L���6~�u�7�a���>�)fk�kT��֡ghgo���% �Bn �E2r�G��;O&e�;V^�z�����w���=yߛK��3�t	����=�/�k��Y@�[���BU �1���جM`����i�.XE�`ܴDz��7�Ϸ��1�Pq�	��{I7��(<����"�	��\�[B.'��֑�Ӊ���{J�����˕�F�P����ub��n��C�z,�Aa�Gt�����g�uz:�h��&	H~\�
0(���o�0�9`2�h�����@���l�� ���G ��b��`̎�[!J���߅/��Rϻ�}��H���j�R�X%�9�1<�����jLO%y��C�i=����uA��-���C%=����F�ת�U��Z��E��Qq$������-]�Ҷi�X燶�c�����"!�.�����G�
A�V�a�r���k��]�C�>���^S�g����s��^�(s:�a�OI�^�KT]M\8�cn�S�I����jD�f(g��S���Z�ף٨��sv������k=�KBxSu��T���|,D��FXU������^e�9��6�Ix����/L�1g���ꍢMa�0�T�X�v���T1��e�k���?涍�:�9҂fX�Yx_�u�9�^�)��͵��C�
X��/�l�ϷH�gG�YP���+�[Zy���A���iT�����⃶5S�<��̷T���qB�_����K
�x��F������ ��oʁ\2�?w����0��r~D�j�6OZL�J��r$5����7!g���/"\�g��1G���f��*���c�z�Rh��fO5���ҁb,f�>M���ΉM9H�W<Du{�1-g�W���Q���K�ie*���FFZ��Ӂ���E��+Uw5�p������s�������܇,����Cv�T^8\i>AP�������U� 8��Mt�D�]G$��X4Z�q�1LU�c5I��Y$2��m#6�a�3�襭	]=�K�I�5e#�����b�]��^�)\t�ф��g�ɛ1U/�`�|JpӤ +���e�+�g|^���?$���`�����"P��.K�P(�A��E|[��B4-��H��@���BjD@�X(���"������[7�dYe����))n���2���Yv��t=��0,5$��ވ�fu�@膓�3���	!E5�K��c�r{<Lb5����b=��	u ���JɜhA���ʦ
?���.��~�w&�&�������E����;%q���KFn�Eɢ�ə�޾�I����Z��Pl_�y����R��盖�_L�@��,��0��x6*m���( v�W�S&oMLWܔ�y7-�|�������F����b�
qA)5<�����f�i�(B|_��nvN]w-L&
���I�ȫ��=�����Q��3�� �u�QI�z�&�>TxO����n��RߟȐ�J��p?���w%F![hP�] �J�$*���n����h�:s>�$����B��L^������0���V�y�b?C;�s�8e�悎ԏ�4.l�C{��q��c��Y07����?���0�UھA����a�
���[����ݧW�B�g���Z����~b)��"��藠�T,�VLl��V'���[snx�I�zy�N��_X,�<�@��37A��T���4�g&Ϳ�Qp���f*웢��&��WBR?${cF�R9*�i�g�IW��8L�E,�oTط���D����7J��ݎ�� �v7�f� �ɨ��G|e�&5�0	�6��y��h�$�^\�l[��e�|x���G:���-�>{Xp�,��f�&A4l+�h��.�F���+JL��j	��t#�G����0�&ӷ�0l���w��=��k
}i�����2
`� �^t`�婘p�t���K���cF�S�10�E�����3Y�4m��W�%�$hf<�!&�	���Pz�V��ֈK�'��x�X�O�z���D� �4*��>ӫ�ˇX߷���O�"�*_I&�����
����z-s(��d5�I�;%б&��N��~X�װ��@i�r�F{G東�vdI(�˝C��_�:��e�DH�r.kɸ̽��g����H���Wmw���"A�K���q?���}��V`�t�<���Q��+���~Y�J-Sؤ�P�<%�]��m�ղ�hg�y�� ����Ȥ5�����Ev��ʊD�`G���N�T��9���������&\�)��M��-On�;��`I�+��t��m3�q2q�x���S�e�s�˷GSȾd´��79�+<
5C�_�����+���A�MĭXmm����h�dV ��HS�<��S9rw�

�%�4���VR����{����1;<ݘ���ѩhB$!�"V��v�I�~�'��4B۴��t���q� ���BI�V����U�`{{�&	�Y'p���s39��Iqf<�A��`yW��8]�qC�#���,�C7tݶ�F_7�:hU���,�k����̩��f�`:�@,�6�G�18k':�����6}�;0����*�Ez�b(�=d�L	��=P�^���A��t����N��~�܃uaF������*ݬ��V��]A6ޏz�W�j�O}��æ���WA�R_eE��Y-����H���G�_�IO�� N��Qg� ]�F����6i��hp����
��t�uP%�N��L 0(c(���;���(�.� �y�Oا�.Tnu7f&* =����Q� �$��ߏ�������y"@-�./QW�j��匷���̈����&���U�M,�	g�AِI��3�;
-�q_��WS��d���(�W�P���6ޖz���+Bu�	|K�G^:{�W��_�#�xH��əZ�t��>�}�I��"!��P;xm�w���#�Q|q����1��Ŝ_�q��`0��x��E�W�-VK���3h٪WV��U������ K��-7F�2`�x�G=�"9��_k����h[$�Eڠ5+�z�I��4�@[� �J�GHI��y��q����졪ҿ���_h��Jв�f1Y���;I�:_pf�W���m{C� ���d��@zr	�38� ��
���#��ff�?���4هp�.&����>2�P��yk�i�^�؄ 1װ�ةb拱�HOu̩��9�� \��wݍ���>u h3֔�trk�Ԧ���P�g��wXrdj���<g]�2��0d��Ҝ��	�$pK,_e��HͿ���>��qU="*w^V,��/8O]�ې���;=� 1�gU�6���}q�̘qjC��y�K��1fL��I��G�g9�'�%T�!���F	�����yDbo�%�X�$>�[E!���<�����BL��}�tţ^ީ?���ȏ��U�ڔB�q�F�Uv;�̡�����H�)�L#>{ ��B�*���F�M���I�f� �sylU��,�mhɜ�U
)��Ǭ5x��S=������̞|�#5.l�P������TO)�B��&�b̤`��cmvo�,;\R��e��K?(�է��o��"�Vl�Ow���H�WS5��]�ԫ28jP9L��־���6���� �딄O}�A�\�����:��a�ƪx�2�{P����ڜ��-�="��ǯ7G���!�)3��/�����&Pa�\���0F�`��q�W9&e��������]�kq"���z���ݢqyy��e�ȠV�U$?���_��Jǻ�������t�듃��](�g<en�؄ AL�w�L#�S��FCi�u� �:��-�IZ�}�<��S덆�;�
v��"��y�?b�D�HN0}Y�Wl�X��J�AK(�� �kx���5Y��%�%�l�A���q�T��o�r�%DTw�V0 ��&�r{K� �5)֍v��)���/�.�4�Oʨ��&�k-oO�T���Ni8Ϋ�N��6@�3�V����i�73�i������0�B�f�HFe�\�@Gҿ����)�	�q"C�o�t���	�~?@�ϟu�֦z��{(>Y�*E�������j�����~5�*�uQZ��ʳ�R�Wg����l��U���������g?�/ӑ�7�:��-�M�C�T�����ϥ4��g<�G��rE&��;E�����{�0�gF�k֜��u�Hg�`�d����)�qQ"��MbV�'³)�k�D�	�P���;z�m��r��k��,F[4|kY��Fǻ��o`�U:��Gni�0W��D�*	�ͷ���'�o��4��维���N���bM�A�X�����M��qh�?�H�����.6�N�wΤ�D����7����ܦ�Z$�rp�UQ�V-˲�۹�H�2q��7��Τ,�ƁMb�"|�����FEj����T��W|>�C�ʄ�����bʋ�b,uŧo�h��.VOڦ���P�fK�����^�)��3�����u�����|��)�ζ�̢�>f�䚊O �0�&e�SC\��z9��
9�w_�]��o��Vs@�-��b��H�_W�����և���I_ϞMe�;;S�"��t��=�mg*c%���eJ�i^�h�}�`2���!w�\�y R{=���h�R�EE&�T߰EնH[��ݑtYj��:�#O[��Kg��ڬ�\�����J-~<�<��܆U����xvc��yY ��߽T�y^�"MGjN���?)}�C�z������4۶x�YI ��� ~^ơ�Fp$��N?�>f_x�� �Q�â�-mI%�[M3���P�1*|,RIC��8�)��M�9�{)+UCn�;��|�^���$�����^B���"�T�F�C�.MZ�A��=|�3ku͡g�m�fcNU~kƖg}�$�%%�>^�
M��TYߊ�SqEB���!��B�{�'�C�����TOp�����	%Y׳��kȊ|��~e���Ȳ�r��q�W#&w���v����|P0ԁ��4�k�����<����_B��u��=�(��-�r=����Y}x�K�{��I���.}Z	%D[��<�����B�z����ڇ#Q�u@��1c�3��T6��~*���g���њ��ȽY*�� =tY�pe��Š!��s�z2��B&x��<��{q��MZ:6׽p
��C�����4N�׆�)ƍ����F ��ۡ�T3>ZA��O�����!�[9�#&�b���p��ދO	)>����U�j��9n[�iCv��B�%'����Z9+jT)Zߣe�I�SX7����[x%�7���9�S�S��k�El���A>��O����"�/9;%yx)+5>�*B(V�;�2�և���Ss�p�A%�t�j:�ԋ�6/m.�}�=�9d��C��(?�G�3J���"�~Q܋���
$z&n9l=�ʝ)�W���n/~�i�Q�M0ր������	J��u�$[�:#'��$I��*>Į�|��=h���lȬ&i U��V%�UU���X�X���d��x���ѓ�s3	�8��K>ߛb5Y��޷�M �v�}'8ZM�T�I�1L�I��Pr��,��:�6i�7�i7sO�=�X��f�����f�e#��a��0�5��#Q�"�z��	$O��Lm��+�����G���;�?�),�AJ���(M�yĔ�a����w���M�G��6�n��L����֠��I��/��O���W�2�4�!�龷{�����GyO)�X�vpv;�O�^�m��ʷ
 5���~ ���`'�����+�����[Y�E��^�����f�5Q��ߡ��q���\���s�F*ك�y�(�EXCgc��Z�ΆSy�w�U\j�Q�)��EI!.Ao�Z�7̱1�w�Γ�Pؐ�X5��-����[����kű���Þ�s��
ڑ���� 6���l���l�@7�M��Z�i��Xr�ag�8��r'֯���)W����Vt�R��j�$���D�,Cu]|b�z�%�J���Tf���6�40%�'<� �M:qF��(�k^��rGM���uL�-g+�W(��Q7x"�L���,(���j �}��X�`������zV����"�G^��?����(�Ui�;@���	�`?�^�G��2�r.0�w=�~�y7~�@++�V�R��y�Y$�����gGv���`Pڪ10y������B��l���ODEX����#��X3JM7p��m)S��VF�L�V}�N��c�a��(��hXk`z�a�4�mpn��N�ILU��Y�Ȁ�nά��[�#�~��z�;������I��ؑR�t�3�^)E|��9�⥀��2���b<-ъ�;�<��4������M�u�RH���b�����B����c���Ę+'�)�վ9<#/����z�:[�|��3�:0(~��\֫G���ᛟ3�Fdef^�z�����k9����X����R�P��fԻ��6���7�����Gb�q(:����hi��`�h��j<��DW��H��iA��Н0�@�wt�s�)�n_8^a�A�&�o1Ø�`ԑ@���\]�F3�)��JmO�lmFgX �ˑ���8bp3s���E����NMl��A/����F�'у�C�"��z7Um�wf�;�=�)��H�;;�&��	��e��T��N��+�yN�Fɋ�p��L��ǜ���zC�!�BA�1ȵGsm-�B?�k�v���Hޒ�Q�"_�J5�uc��*Y�x�����j6NX'��tM��z��7��N�2��D��~ Z�B�$�7�Ba�:���|Չ(-��>I�;�F�}���W�B�gc���P]����^|jq�v�'��n�F')(w�B!�yI���1���"�([�8f�����3+��\�M��A�;�&v68�%��2r��|���ԗ-�3������)��d g$�C�b~���-���>2��u�3�a%�K��-�L<��J�Y-l\ֲ�]/�̠��k��^#��'�x���A���.�I�En�v٠M�qB���s�&>p�r��uܱ�EV���k��-�q�0��K`���l�ɜ#S#����FxG	^��=�*i�By�t#ʤm�1f$D�t���p���#Dܯ�8�?�)�z����Xh�;�_����pw̴G<,u��o�l�"L���e�58�.�5l�F�(�����8+��Ҙ�>�g�+%�3����T80�m���xm��n�A	�*�]�+�	�u5�=��}w�]�oޱ�rtn�Ȣ���`�|�H����[�K(5S?��j���#/,>�	,�)|-���Y��J�[9v'`T���3I-�w��k��eM����	��d��EK`,�������8k_.)F�-~W��Nܔ���c������Ӎ��O��R�Ƌ��.���"��\UƐ�o�S���H��'�[J!�S���UR}��a1�r�QNV�8��l�N�����HσH�!��}=�b��'�̘P�c�K����4��F0��E@N0�W8h��z���'�A? �=Fԫj5�F������܊�F��� �8Ϭ=p`�% ~�Uv�\�h�0F�c��r�C�[��?��	vT�bƷ��Ȉ ��=%��_.����¦�	N�������۳�����UDC�iۀ
��vlÈ��OX"�ӽP���v���ln��.�#�4 H�8�j��7�z�w�:)v?��Y�*�ؖP:��)��t$WR�9�!����Ƣ�:�����rV�B�ɚyE���q��xƯ���Eק�䟷^���HL����h��H��1f�ϗ�$wRvd9~X�-y B"p��OJG�'���0�K�@M������� �@��Ǆ�qf ai���'ȲbX��l���_����,^����+���+|��XjԹԣ����RN<�g�w�;}��Cgc�6W�*��"fc�����H��{5�ı�F7i>�-��$���my����bLu%
���D�-�:��2��%~55���皿���[H�|J��6�\��u03�d���	��S?��[=-�����<�)/�x�})#�_|��b��<��W2��8"���ps��d�Uo�x�����yR<����y������R��U��>�mF���}!��o�k\f��+�Aj���S�+r��'�3&�"��3��굛ׂ�[��0�dz{V�������ɻ���3���?��~Q�I(����kmw�����//�TX��ʀ-�Zmr��=ՠ�U�YT�z��䴤�|a���-7��q46[l\,�
��y���B�lj��I����H>cY �n�*��{w��Z��ժ�޹��BSZ;^k�|v��,�P;�*)�~Q9J�l�^�Wu)҆Jʹ���L���3����E1�ً���"dX���'K��/�YY3R��N�6��$	���7�\s��V$�Y���S��j8�:.�Jw;D�BQ��!R#�Y��$�����;W�@{��D�[����[8�k���A��?��4ȨP��k�VnK�&CH!l1h��"�	�`�P+.�,k�=�(��C��\�	�O�f�?dӕ6F�v_��H=݃�ݒE⇬�sx��6;Ǡ�XX��$�<�C	@��-���{�󴄍8�#x��j����эșMyő�jL��k�ᬶԙ�& �m?_��ɪ�y�l�|��ӼF_�#0
���ewF"6�?W�a�S�n�w �����`e�5!0�m�[��=�2)��Y�o���s]��g�༡c���#b�9��:9q�H��1Br���Z�R�фv^��=�ˡ���Q��S��T�R����H���h憷%���y��b𵫋��Tq�3߯t~(��I�2���#�z;� eR\��$�����r���ٌ�� .����⽛�?}�W�l��k�]�"޻��A'/��"lB�١�b���#�鴵��dU�?P��yx�'r;�|8_��{UKL�(��j�� 8���왋�T=��9i(��Q��<��(a���tY&6�D�Ep?p�5�2!�m��>����Ȣ����K?.y��z5*�S��9\�yAg�m��sǹet��q�E�L�jxدX;���4$h�ݬ`tY:��r�?�LrW�=%P��ǯ�Ke7��)>ͺѦ��l>s�h���N���"g�۝"�n.ZR4�-d��n���n�.�E��� -����cÝ3/qM�XJ���"�A�Q^��7���������I�8׽zN9��ٷۉ��3�o���#�ŲG��g�X%��
�"	M���9��6�s�����T�+�t]x���~=��d5J�@�c�%��[�O��Dݒ�()y�Q]8
�?!��������d�b_��F"�z����N��6��w�m��&�C#�|N��M�Wx��A�H�FL��
���jm��)o����ݯ��(����EΏ�%E�ޕ��bvzW������f4�w����.;��gA0;�&�Gics|��{�*߳�8E�[f-ml�bsͦ��������f+��Q��{�gQt�]�9��h�i�(Ev'����=��^\X�}�P Kzx�;*`�E�8<�}�B�،�z+��_U
��w6�9]Y��⨤{�#7�B%��(��sAP�my&��K#�4��w9���y��b>�$'�2��&�K̖i�D��1b�k�z���;��rEyH��~?�t���5d�]�ǇW_�0�#'�b��)�kY�-�;�vɞ�밦_d���8����Wo�<ܥϤ�@O�8���ٯw�Ҥހ��r����:桁��Y �����$G?���k�RC�_R؎�B^j��?\X�-Ӫxl�(B`�����g�Y-֎`40-}�[�ݓ[a�o���m�JZ��r�3=y�.1R��������4!�0��>F�7�WVt�W��Th���\���1"��������I�}���S2ceE�/��1���,����?�p�8��w�C�&�-�m^n`O�\���Ńs�#)���̦�JQk�:P��B��4h�HED�+�%=�%�2!l���C|rvH��G����7M�|9�}g fE-g�?�w:ѱw�����(�b�&���0-��_5�K�"��8��h�p��N�+P`�mWjA�լV��		?�V���+�L3ػCo�ʮ��U�����,
�E�I�(�mm!��-S�0^��#���R����t]��IM�N�5u�I�+��_H�C�-��G� ��<@<(�d�����	�̶ѹ��Ɯ�uy��p$��n|�ܙ-�B���˟5D�96�j��7O���_��C�<��i��m�s�5Y�2�������̰�ʷ��ö��U�E���>�ܖY�d��B�)f�{���䝨vD/��UG��u�6�~�)�����
�5�߬1�?P��{P�"]�����f}�4]���b���K����7S����b .D�#�.�/m�T'E�wl���/y�}�~�5.����!n7�I�A���r⺎�y�#6R�}I0 �cW!Jߠ�z�z�F$GK=l�r�J���ux���q+�5w@�m9 ����A��P)�����!K�N;uqPh]R��;�㾐�%]zZk�|	��^�,tCQTxLn �Ɣ.���}!��
w�l�mP�ت��(Yߣ&/v;{����K]��`��FZǃ��:Y���3��e�rxȌ�$����͓������Si�SJ��b�5�����o� ���_w��Z1�lP�V�[*�i2Q_�x�����3O�Ku8�����R��V��u����!�\���%�c�� �hsޗ��ߚ�� @>G�&Ie�W�A��o_���,(	_l����`��Dy��>�\m��|ޥ��f��b���Q���m`1t3�$���}D�k�x�t�e�E���$��o�l�owoR6�)yۭ�O�(	%6	�Z��Y��pje������)T�B։H���"{�n�fg���(=u<X�����<y2�n]���w�Ն�V6	�./�����YH�9'A���\�ձ
5e2&���N��o�.���_���#%jd�583��x�b����83��A�_�-�7,��Z�e���@w�)���X��%����Rv�c���/M�m�!|?��&�Y���sZnLR� ��ڒU�tY�)�Vx�`eɖ9r͝{� 7��A��;]���Bjv��X�5�*��U�y��nu�nߍ��� �����9&/H4�"&��w�O�`"!�R���n�t�yc����Jfl�y�/��R��z��^r����_�2j��9?�O�*#�eFO��5}N���D����V�MMX�~=L��d��6���L������/�K�`-b�ue#`��% ��I?8Җ���gv��e�����7�\�y�$b��J�c�Jy�ĵ
�1��Pu�}�H�dǆ�Dny�$@ҕO��5l�^��n�;k�	W���`_��d��;�Y�!�K^��\�rD�Fc��mژ�fS���M;eJ�{���?{���M�A��J��ƥ)lw���ꜿ�E(���!}�pM<T�iUj��ʸ�����Y��v��m�3�h��}��F)&x�q��<9��ƦT������e�Z�(�hb~%)X��=���
�&Y�%J��v�����WK��<+I��X$N�N�15�H�]���%�\Bڽ6Q���c㳂�3]`����x�R�����Y�Z��n�r�x��X)PX6��/3�c��/�U���P�6���#����4���iY>���U�r�S�956^�1�L��<W�����.���X��:] �����f3F���� �0TB��c�����P�z�s�R�$�fP}�HNY-] �f�(~U��r�jׅ�` �,G�J��\1���}�03'{��2 4y����K��(u�t9��vD��k��` �W�p�կ��M�y���ȱ;˻:�͉�S+�� c^�y�ū�~׬I�L�7d"P���jm�K�^�'҄��±Z��_r�a�O���iH�����T����3Y��52��@:�����u�27o"-�҇m���b�%���{�1���o$cF���(���s�����:�ra|����k��~)(C�G�<Mq�3j�Olŗ��1���ʞh��*�|+K#>~�Qq�����˥w��z��/����;"�O��<�eI	R��G:���Q6���E��!�1�^�Xxs7�@�4[�h�Ө�ĻT���?�E<���=Ffe[�￲��(���U�����vcs�gbP���"���L�n�F��(k�A����K��G�3�ݙ:�~��\��:�s�|���y�<����#�i�/)گ�ǿ��^UR��@��pc�#YIa�PL����jΡu�?�i�N���b����T��HFu�kR���J�y�Wl�m��/Ɛ�Z����\�'�X��}ŖY��=	`��H�r��RCIːsP�)�ſ"�>��1�tk"ɳCc�5$ ��e;g�o|�lgԱM^6d z�2>�U)�=��u��u��8�w������̄u~�;��`F]���&�!x�lExKĄ���M��!~)�׉�]���|�,��b(�i���m�b����,d�n��4F�vD�� n����OE�=$�movH�B�,�{��k̖�ޭ�:�ˡŸ�,��J鐭�T���'���ۂi��r��@a�[3����0r���S�F����:,�T��d�C~��?�.}��u3��L%�q�l�>�ŀ��%�mɽ�x�f�]�\���Ǩ[rW0�?�>�)V\�>������&��3��f]��W)�r��4�����e_N�>��[q�� �����M*��AcvkCN�MH�M��_��7����殛�G6%$+U�S炏*e#W��7/��wdg�&m}���u�d"��܄�5��nĮ���q��1�����O����y3�W[X��(ꋇ����;�N�m���`=f���y�Us&��H���88c�Խ��i�>ADYe.;�l��"���`"m���q�(u��y�<[ڴޢ��9��f�AFGN�N$�i�џE�w�1�#i�'[��� �4�iJ�W$��	x艞��R�ؼՅ;pn�Q�1��_���Ѹ���=%�
/����}\��o�����}�(Ft�n �E�:���§E.�����t��*M�e���	��Ϸ����/��7k���ч&m��c0�P�p��R�#�7��y%�u�̎�ߵ���[���0%~������
r���v���h�v1��>o�=Tڨ�/q=�Ґ秒�zOh��q��r�?�d�#�����g�����:�`�gs9Vn�ĕ�������E�Кv�k�a6G�Η�]O4(���Lb"c)�L}{Ѥ~��GT�E���z/,��-	}h�g��igM'�]�o���_A�q-Lգ��#7	[h�U�UuQ�[q�4O@@���sB�;��N񫡒�Ĭ��Q�=��BMWl������9{�1��n�7�Я���Wڡ'����H	�^U��ق&��@V�v%�>J�>�ᦅ�������m���
�5�#J�"�X*�&]�u���	e�m?*wʪ��{َ�u�V�ޠ�DiR[�3Y��?�bE��,UB��a-`�e�\�n�p�	[p���r%���>	x޼����7��Q~K#缥�<�3"�A:e��U�����g�R����Ҧ��H�U�I|�6p��� L瑽�m7�BI�C}&;%�zkY�;��V���y��o��Sؖ��+�� ��b���L�f!iΊ]-.+�H�2��ĺf2��`��J]{������ڽً��e��r��������4�?�Hd�����%zz[Y���o?B�WJڷ����jc������V�:�g�hb��I=��4֋8̞E�	��JR��v�ő�Ǖ���N���]>��<�Bh�~I����U̙^��%�?��Y	�T�F?ߕ�h��Uu�7n� @�:�)]FWM����4h���b�aQ�>a�e��ڃ�M#$���f;�5�ZȜ�z�~NjO8?o��n�o}���_��2����W,M�21o1�ʉ`��D�@p3�Ƹ�qU��Xҟ�D��.����^HL

�-���@
4<�Z��V��Ǿ�&z�� G�5X����)�t����t���7�$r�����r�t�
�C�_ML�Gԑ�*
��.Z��JT:gX*<�#�홆�u���>�I�H��F.���y��Li˿b���Pl<ޘ��h�&q��w��41��T��2��﬏H./���ȝiTt�������K�a��<]�ivn����x�dK�}���\im�\Y��&��j>�J׽��Mo���*ng+>&�8pO ��l�I�?�%�r������U�
U,�y�ת���v�V����J���G^�;��8�r���"�i"F�FV�1��?	�7��'�:xb�0�g!s ��&'�.��i]]��W7�˻q6Epm�)��7���9��p*FQ(���6RUE�dГf���>a�0sS�o�y�H�+�l¶z� �x�<!�}���#$���}F�NP���_�����j�v�͜ٱ.AhW�Cr<�nB�H7�":H&
�[���%9�S���ioJN�D�.gx��X�G4��ZQ�z�m���AX�����/��K��Piw�e��˧�C���S�5 �썫���]A�"���e�цeܿ��qGfD�ꠚD�.1�戺�lB	y�i������+6ݞ����D�
_z��6GM���.����˶�LTF�<��9������"3� �o�֒߹�5�J��o���G����e��6�Y��p�)�t?f
G�h�ixF�U�2}$*t��-�1��p���	����j|�ɧk��:$��+�E�!H�����*@�*m�iԚ	3I��j���9r��1�Of�K�*B@��n�\�7�� &[V��5s"����ǥ���vx5=e|���1L~u
a�g�S�i�1ɾm�m�������n�Od�������MA�y�9fIK�o����՝»t��)���.���sX(Ya��*
IJD�*HrՕ}�׈�y�gM�~���[o���?���JY������ef�[�g�����Ѕz��,��ɫ���3�v�v����ԖZ.Y�C��@d�hR��˄11%щ����5}��.�=M%OQӴ?ÿ�Q��yȄ^�(iޯ�Z~ވ%�#.Y�Dɝh�X6�	�Su8F��C~�5%|o�"Gi���1�(��Y������V���p�e@09��y�� �x;�0�R�?M,�ϸ��T0`4:W�O�S6���9�>�ݺ�\�g�������EH�+ak�3����+�"��?���̰�hr|
��磹�i���I��������B97G�0���c��X:�v=�PUk�E�H�����O �f���z�� �����/���<��� 6���x='t$�xf�2�6Ts�_$xp��$���NW�gێh�E���R���'J�BC<Q"_;�e����&��Cy:
@G�����〷�%�in��쾰��9�M3�~���[���(�.~�>�Z��U�o~: �0/z&_�P�gV��XοHųTE�:t}��ٍ�?�'�c겞����C�n�{}�IIS�����ű�!���8��+��ߛz[6��0���ӧ�?i���u���L8�oE(��r�
AhO��t��{Sf������p��@�r"œ
�)�4�Hx�%��8�P��w�[��Y*����j�7v�	�p0�_�ʪz=����$Ǒ���
窫u9R�D&��\T��bd��ߩ.�x5��	�$N9{�}�� � X�a�4:��T�u�.#vV�hX�u������{]Z!�Q��z������&,�!���+�\cg4V�L��x)�7���T��3⌈���Bp0F�*��p���"F�)U$��H!�n����[-� ��K]g��Lt��V�F�'ܜ�� �&�o��p��s���]������"j�IcP�0[$I: ���[#;����V�KȐp�C�䀈d��UnH��δ�D{S�=qZ�Uk��\m����R�G����m��Zd�? �}�/z������{9��r+
�r������Gp[~<Zʛ��e^10��Ϲ=���zx�M�J6���[�a=	��ҷ�t�rp��K�î-	~#����c@[�^2��Qc���x2�mi�8̫��WAc����x�ל�B���#ib2�E�d�:��9�{�a�W��������	'8~>@�eSX�ٌK�ʖe�L�h��vK��v�Nz�f�݈O�l/z	f�v��Zߔ�:)X���H�E���e��ڋ:����`v�Y�7;�)�`��t��-�`]7�� �%+*Ұ���嘺����?�����E��< �nu6? vι1�������Sd��*����e^G}j��a�c\��L����q�a49�e�����`�<��.�L-辽 �~��FF���k���;�u�0�S<?Z6��^}��'�$��
�m{`
�{���W(�� <K��ť�39P����<�Y=��7�M�/Q������7n�N�i	� x����v:�s�!Y���QO�V�f��"�vu�n��{����e�@��I� �*iY6��C�
�A�l� �B�;4%�˭�<<?V���ǥ������w����+��p�]���?6Χ�߅����t�1|���V}�Oo�(RbW� Us�W=��7v�zb�C�'���:�)ر�I/��f���'Ŗ:�I�F솟ϵ>Щ��Z��d�:���:�\�$t�Bx��?��Z�	Ӥ��A2�Iݝ��O�;�oݦ*	WV��k�2�*)TP�90(�f��<���آ�;դ�Q��֭;*�K<:L�+ة�����2�Ҿ:=�s!���r�b򬈳�������>r�x��\sw�W(d0�p�?Ǎ��I��z��q�z�#*#ۆ��kԫ>��N�6kN�R�O�nҵ%���`�J��mҹ��K�%.%�[&�s:w(��lv���K��d9
�J��NT����?@`Ҧ#h�ёs��b�5�H�r'�1
�o�p��6 ���A�bB���n|\X�-�ux�2�=��}�ě���F�0�rO���<%t�>�;��q����Tɲa�a�tЧ�&�.cw�+�w15�� U]�w�D�l�p5�M�d:}�d:R�'��=�����Ѿ@�.�%D�o��"�f�$Zl��Ľ��r�16��Z��&�U�Qq�?r�U����t�w��5Ѷ�� 0{�2�~$?�����K�B/��w����+�`�<����Ȫ��A&�K9��A����Z1�9�B4RH��RZq�5\8w�*�ߗ�Ok�+�/o@�F��ҹ�gVy����N�2�����R�5?��D�XbD��؄8ިR2�o:?\�{̑JgMӭb.�ב9�$t�6�=rɶ�L�/����{c��t-B��kCֈ{�B��Jg;�NA�|�D��Ϊ묪��E� 7`�*-�Z�  �čn�ˬ�� ���k�����Ã�?�_��$�j蚍��kP�~�^}78@⅀�����m_�a��?�K�� ��Aǁ� _�&�2�Gdm�qqxu&���F)�H�3�Q��aՄf7g�{q�/B)wZ�i�c��L8��<u���-F�[x�8����;�Y���R����,֌�Q�84��C0���-�6(�=�E ��K�*�ѯ���s>K{Z*��d�yZ8�dM�2��Ut�G8�9$�����jd��&�_Xg����uh��ß��79ASF�]�RBx��� ��X��=q��c��>m�! F��
� 2e�{�q�I�X�Ԙk_���ܦ����'nz��g���7:�`��S*�K(���3$�ȬM�O��C�ьs	��I����A�՘:v�xtt�����Q Ε�_H,�L����^��5D-�#¼k��i ���{�C'yE�[��m4�G(��[~�eA����@}�h����@I��ϫV�P�J��q���ݭ�. ��&��<Q�>u��ċ-�En(��?�/�:� O�4XD��u�k�x�	�dJ��\*uT$N5v��ؾ�l�7[�	T")<B�}�i���U0,%e�W K��OFO��A�|PAY5��|�UŦ'h7�,�.��9i������P���˾��j`�u�)�(F��<ܘ¯gٿ�Qj�c��|������n���<}1���p�
=�[M����c�����c����K]�D��T%1{��!%��s�_z�8#�C�cߒ�=
�-���T��n�Ș��C��/%�q�фO�פϤs���ō�2�<k�A@o'���|�8�Dč�g"vZ~'}��O�cح5;�'����- ,
4��Ȳ.~�~������w��/d�8�?��������]gˉΖkWj)��Ix�r�72�c0�M�$J�c���.=�c'���٥d;v�)xj�$��z!�F(:�Bw�v�h
}q�c�{����_�&��Ǣ�60��Sּ�/�P1G`�z	:�+nY�����
M�@f�Z�E�v^�-��R�RT�)tlW�K�,E��C8���ו�D���4��W��r����1=�z��Һ�?9��nk`\�&t�B�Rc�)MC�rJ*%�<�?����Ԉ��mv���?���ܗ4����w�G�c`մEe��*��>I�<.��2���&��(�xt�Xm��
�w$�	��D���V{�-�suT���H��*lZ�1�H g�N1���m��n� y�ø
�/I��е�Mg	P<>���I`��)In��s��"w��x�[f�Ƙ���h��KC�5�jp���m��1(�#;
Z4���	o;F��p����j�L>L��²�Y.�T�iA���8�Y�<)�����$t��£%�:RTъ>�d�=���*RJS�(�j1A�P�Abªs`jo��4�t���Jhٍ�|h�"�L��� CDI(��?w�^���(]�?��LP�J�X�� ��܃/�$��?���b/���9�.zފ���Qk�%'�b��L��흎�?38`d���%(���(4w1_hf���i&�27Uz�3C'�M��Eì����C6�)�MG�̆��=|B9�����������͘W/���^5� ���?��b�R�;����۔_iY�-R�&a�"Ԯ&a*ݯ�Q}�V�/�y �J_�L&(<0�/r�����(b�wßҽ0�yf�.BY1�I,T9~Ya�,Ge�L%���"2����j	t��
����g��K��Hn�|I���ڇ�ųv�D�M���(R�xp�9������E�I}��c�����8f"(�&��k�k=������2�W����b���拡���k�{�ڎ�$hu9�vq?���|��/�'���]eH2àH�0q�<�@zYE�@/ݙ'���sI�{ L�%�lD�e8V��$����� %�r�k�%��Ǵ���ՙ������̧"��&_�<���l�m|��`M��z�������Y��\����js�6�?��뾍�Ϗm@�ma��Լ\�Op�㒺'���׉,�/��x
�� <\3Kv~k��9����Ö
3�E�RJ��(e���(0Q�mI'n�Y��}G��F�yJ�JWw/w���Zh���3F�o+���n� �A�bK*���[N'm��7������,�t������7�t�h��Y����#�&}�*�8�1�v���,W�:c8����=,���u�k ɞ<B�eov�����Q�@z�5�N"q�`�0�r��9��LH{X��n�gYS}GW�~�ɦ@��,�	'����X����ks��4��HEm��M���L�&�{��B�	��]���� �`����k�ZhuT��:f�۹Y?q�p�������ּT����[F(���r���!�q�nc��վ��u��~ׯ/��=�c�do{�"���]�����{�܈�a�xd?\�hRP⺢[�t��s�|X��$��Y��pˑ�M_�Ճ�T�ofջXkH�qV�����K鹥��9�tO-����}"#2��(��5;^Su����*T��/��)ɐ���3D�u�Ӳ��Ug��,���b�V�T��U?ύȶ�5�F	���C�r��i���S"�/�ME�������E<��͝*u;K�Aݥ�ɺ]�V�y�<�)�$��0O����]oو��=�5\	�q��x�i�S@��S�V Z�Lbx@j���N�8�����	d��Kj*��^�P��S�{�c8�٩t���<�L��3=���O�? �8�a蚱4@]틕�o|��q7�0=���X��)�}����:�>D�D[�5U�C��z����7���p(����X�p�՗p�J�O�S_]_�����Fh��S�sv�7���O�����;e����E87>	"#���Yۢ���θ�^7��P��Hmb��^�Q�SH����������:�j2��2�M�P����2+�h��$���t���5=���_+�
�I� 3�*�O��Up,�����CǇ�h�Gd�W���x4,ga@B�B�ͣ!�[̆�U�4݊FR$ǧ�pt��>O��b��X܃6]ZL�X�	7;��L$ᷢ��ly�s��¨{	�d���C�� k�ae���죛�}��(�Z�K��&<���Iy�yE5�]$�w�sl91n�#s��
��	n^������J�LRx8�{#�x	Y$$��&� �8� ����T��^������e��0��k�nysP�������j]|���@�I��뻽��7�l�ێ.	Bc	��gj�N ��S:s��� Iw��[!�f� �;�2�P��XB?�D+��9���7Z8�P�ji�C�M��x}��r�3�]��P��홥�@�[��TRU��q><��0��TW�D��!v��.ZW"������F���8��Xj�X ��$����3�)�4If�4�x�Y���DŴ�JTnFB�z���nNW��w�wg�-)��������م�5�*g��# �&�.0?`_���/����k�<{���Lo�u������;���;@M�����\�}�8���E���Oq|gOq]��ac������U����mv��㫃2�4M�d��{��4�,,k�i"�˂�W�/�| �!�t��G��'�h2�,�FY��|5�H2brd_��&�z�F�t�LKU�*1�u\���0��)�|�-�ό91V�g��7P�)���
kB@9;�SFNmq���3%0Y��sMbE�VFnH�g��a���"���q�>�YO6��6��׹�>�`���~7o���ud���e�ʾY.Z����\M_��8H1�S���2�J2�ܥ���K6�:��.���1�'�\Zuq§�h�y2�<H�E�n��0�'��s������up���%���o�=��h��Qgk��-g�?�^>i�y����.��,�Z\�1�����ل�Q9�f��f��,��_�<s|����	���Hc��l�'��������J�)����oo);�I0��K�&G�����H�������M�4%JP1k��7�ŭ2^(���,h����vщj�3܋�x��e���O�4? �7����C��9��6Nۿ�X@�*ѽ�'�Ȉf��?���Mz�Z��`��f���k��ԅ3)I<��DJ��Q���X��y����~�u�9�O�eͭr�S�W)܆q���Cr�`�> ���N�_�&��'�4���u"��&m2u
$c�D�=a uK#��S�p������w^�?L��$,�����-I�tM��[�:O??D�ø���h/=g/k�f;��j���cR*Yu7R[u0�h�Hi_��z豫3XZm��CI3s���{p����ꡰPv�չ������cv�vM���G�7�B�
����gI<��Z���)킡4�-�k�1i���nh�Sw ��
��M���#d��}�T����-4^*磶��dd9�q���{w�y/'.Ua��2�q�(N|�=��Ǜ�Cg��=������<S�i�&e��6��D��I�Wr�]���l�-r���uO;���>���?R��쳐�g��{�~��}v�N�$���4e;��&V���m���SN��i�	x��K^pѪ��p�X�R:@��c�X�D���-�F���E.�/\���fވDQ=�H���,FeI�\wr�΢G�y�^@�����႗�i��Y4狓�Yz��z�N��s2��vX��U(G�a)eߣ�0md�	�>ߧ�|�0�U.i�̠ݭO�70P	&��S�S�<D$0���ͮ��:�ϖR3i��K��Qk���u9����ܤ���߽�h����@�k���igO�6����e�B1��7���X�f�������$68K���n�J�L�U��J�,������X�ݥ�]��5���w�Q��l�*�E7��h1/4Ġ��+���͊�0��[SkY��k�e@���S�H���g3;���Ջ<���ڧ��O���O���k���	޾�/[H��6��`��-f;��l��L�� ^1i�PN�r�'�b\�P���a�f�GP���G	���E���7��K����o'oN��8%�c1=޽Ɵ+> 2k��9��1��N�'����s�[Tj�KLu>c�Jd��|�
����$�٬��~V�֫p��+"
���!��lӗ��W�.U�C�{[�Z����R�爪�/Q΁�U` @�g�ڿi��#-*O��X�bv��8)� [����z���p��l���L��AX��A]�E�����j�h�W4_�OqMU�x�kL3G(ۼr#�~`���:��z�[-��6�S����iFh+w�>�	\oc�C1_����� +n�f}�����X�c�'bf������7X��� ]�xB�w`P�R�̓VM�i�{(qL��C��J3��ӑԾNՅ\�-a�i��P�x  �m�2���Fá�e���E�C�0�;u�X��^�+z�p-tl���1 ;�=��B[U,K���xy�`�g����� v8/�W'�)Y�#��kk$�d嗁����$.��t����`#���V����,��c	�g�*/�.�R��>�KӼN-"V4mc!c�+�&c�ǔ����|�.9�U���koM|����r�2UM��N��n�tԋ�Fz�(� �!z���t���ק�Azr�f-��,;m ����d�&���Y0��R�j��ˉԨ�0��c�w#L)�}��2�B"�-~�I�]��$��'"Ǿ��m���m�+i�O
c++�͡H�D���)��VO�^*��=�e�EY-��[9c�����5���D�	i���B�����~�%K.|jYv�*ᚭ �7*K4�3<&ma"/�W=��+���Rű�ڮC���a
 �h�ս$]�H���B�+>��|��Q��Ҝ��\��~�� ��i.���9��w�.��T�F��W���tx��.%B(D��"X�u��:g��29�uə1K�6���ǥ�#�މ�U��ഔ��d�_]&�{�����6h��)�����	f~�o�[,[񐡹/�;�ם�<9(�!<�V��4�<E�G\1��d.hhOrTo�V�w����)�ԟ$մS�JGJ��ij�����0T�D<�sM12J~�->M���R�YI�w ��j%!��hû��vt�V4ck��MR�akS�L��W���(��p2��jBC���՚���e*�~C��	��։��	�"�	wc5m�)��}�C������K�*w�C��TW�A@����n�ekS��Y�0s\�%G�x?�N�o���.I��-���?T�Ǣ��A�����Y�V�,_���c�7iD�����I}�E���z&��xFBwt�b��W�Y���5-�P)5�7	P�=�ł�q@��Z.�&n~���g�z!�Y��dF�[L�"L���P�FC>��O�L;��u�O�۳Ѓ���b��K�~�����qv��}�""�����0�l�FO�S�������gya�`R���pLL=�Z��Ǩ�D�T��̫�w��P���Fޭ��'�N���f�kiǱh����y>�|�I7�g��'�c����"�����Ʉ��T��G.���K�j�U-�N6
p���/�Vbx�A���3(���IYU)��"�?�xN�\��͟��+�xY����?i!V}���L��t�I�ul�!�	�i�wX���Y�u��VFX*J1���a�;8l�����m�b��\EM�`� ~���t�mUC�
�����.$vp�h�G��:h������r���Y�uB�$Y��	�7�\��d��_.�U�v��IB���mq�h����B��3�_/HB��`��O!Nk�s��l�*�Թ����w\�E�����L�2x��/�6�w�,5P�*-]��H��D�\�Ta&�Zy���j$}O\^c�����:�?����P��\�>��i]�y������i�޷Y��t7�!~� �]�0�Q�dٸ�8|	���:^����:&)�D��W�夳1)�iE���3��Wű��Ry�Զ�8���*(��¡H�a*�K(9F��:�������=6�n��~�`.����{`�qjH�-�[#(��>��I�"��;�K��մ*����T�����n�O�{�v��koD��~��ī>����<��SM���s�F1����n�`~9[�� �]�6�6jw{Ł�>�]�}�]�˳�{�'��w���m/Whg? ���si��o儰�_�9C w¤i
��	E���&��yIЀUk#���ү�>4��X6�aA���o-���a���MIVg�4�&�h�}�ɼ�4dYk*����Jc�ۨN����{r/�4Ď�+�*�!οbw�v����Z�[�\�>�\D%��hԚ����7���u[]Z�8�5���"��H�8�a�������rO��k+�8AZh��@J�i B��py5�Q�]�ԥ��"i����~ɪV�Ƣ�T�� R��kl�p�ӛ�Q�|1��L�M�X��y���ށ7buC�>�|��]	�$���2�O�+�3�YO؀��6�Heȃ��fmV���յZk�M�&K�=�N�1�/,w����J��M	��O�� (Z}lK��6�
���(�9��H��3� �6\<�/��1;�N��K�vG�1�
�>�NE�	-���H�΃�~�0����O���$���Ӟ�;���hy��j��MKn���L"��ui�"������ �Z�Q��7*)@��ʔ� &e�G�t���=���}~���d@�@
�&��i���!��w�G�x����jw��S��{��I�xHj�P+o%f�/^�:# ����a�I���x`�l^zR~k�_����V�u��Q���sS[,&g�d�2�)��ײ*��/�HѸ���g�}�"K��6�j��DAWʆ��x�u�W�����j���y�ʿ�[�:!����j�V��,�䪚�Z�7?��TP���z߰0�ByX���?[�_,ῲ�0?�m��)���>����?�J�l������h�����6�����ϖ"��,�-��߉��fl�B_��agϖ��J���V�8��f���x?�����@��R�_��5�)B���8 �t�V�*�����cӱ��Z`���?|��"W%+�!�����P	������S�!c��]�;�vN=��w�,�ɒ�$��l?>��'E:�W�D�#��%O����3�0�N!I�;a4�ߐv� $���<�Uhx�����x��1&[��ݷ�*+�>���TUmFΡ���s��_�ًk����*@	���J��gCn�Z�	[�����q����׵0+J�%@��w?���{���M���UAF��PXlc����=~�V%��?��D�s�死�a C4�s�]IT�ίD�Υ���xxg���(}Z謴V�H���y�O3�aS؋`4�4�6kg����-\vޒ�z�y�6�52��d��Ʉda�O�2E[��+�K[L"�L��0qc�볤D��\2PO��Q��:Q��������Lv��>��)%c��G#�:�#컥d�Y���[�t� `x��;����M5��ڃ_��<��kvz�1�(���z�-h̡�`<Hs��M��<n2��ߪ �L&@?m�"�\��7��&L���^ϲI��2��9�,-�'�O��������㢟|UXe�m�襡J����PZ�k�c��;���@<o��ꩮ($Z!��N)� [w;�p� m[ӿ�IƆ�[JA�\�I
�ߚ�6�o���}���+�Q�Tο�C]��._��o�w�=ս��WS*��.��u��
����������cb�r�s��tL��
� ہr��㋀�;����A�T�����R�Ǹ����I�f�f\� )�i�
��Jn[���$���b�d�Z�a��\Hp8����P�>}���Z
�]<C;��*wq9ʻ�|�Ty��	��U���A�"��q�s�n��4����W�{g[DOW�R&�2�Y��)��� CN�	�\*Mv��u�P쯬u��	h��9��U_@�N�3=B���.O����.- >�ϣ6##k�9�;�� ;D��oy��y�9yՀ��5�aƲۿ�� �j��}t��L���D�D�p�}[o�/ϊJ*����>X=w.<G>M�D�0�[YCV�e�0����=�e�u���&�9���]�7"!lȅ��)�w�Q���BD2Լi~�w'��my���\�K!�7L�ƿ���������B��d!n`xN�c�-����9���ൗ�Bbfe�><�*� ?�>_��ޡ7I�a/�XE���(ː�m��ܭۨ�Oӎ���9��m�*�4nQ�	*�RNl>��ۏ� 1����"�	�������r`��K��&/�Ԥ��2ǯl�*�����M&��pM���.�$�4�@*�@��uLI� ���F�4��0&`���*(r�\'lK�hab=�\)Z>e�kY��bM5�y��ܳ@N��^��<D������������x� T�_�$��^�;�~5��"�{q�Qj�GVx�<�]J�凬Ф���k|l�ޮs�i�[&fn�~���!f��d�	c!	��~��f��������@m� U�tP{�� öV�oR�u��U�ſǺ�w��lp ?��B����2�ww�G_[����]R@I��Q��^.R&'�u~�!*>��α�kVFO~�./��Tf�h��׽L8ߊ'N���w�׉���f��
���y'�'er"�P��Ͳ��Z2k^��=8m���;�2 �:J�]�˗�/mW��$R�ZkO21���B/���!Q���?i�Ng��4Rh��ke�b"��Y�l�O�{��N�4�`�x]�> !�aVrVSyp��m��^�ɸҏ�g��F3�0J��_6�@˗z��d
sa��KhXW"��W[Ԡ���83n�w�1U�)H�������\�w��T)�G���R��WZIt #9G'�cn�+�r9fm�g�+��B,��9��n�G�k�Ef�I4���-�=�֒	8&>U�XQeg��!,^}&⍠�+=�X���DU���e�Q��ܖ��~<G���u��A��<~�5��C��`�Q�Z� �ӓ��휕2ʤ���{�DO�uiu�j�5���޿�͝]]�"�AvePt��M_�>__Q���8��p���2�X��"Sb34�dU{��w��|�"K�	GC3�%x`s��t�A��ں�~��~�w�fU�n�;,˩v��Ϸ��Ȫw�o���:�S��W��fGȿ�� o���� ����ѹ�'�嬕n;���E�u�(�x9�˻C�-�SǍ�� %�	�ȹ�����)>�U�H�I�����%L�a4��-3V�ʗ˹�hU#�^��
��1�i/�����n�O>N�� EK��d���c[۲y�ð~v�rV���b�eh7�8��X}���k�V���}�ٛfxe���z��:'���I��o+��UX�@��~��P��3-�3���4�c�	S����wF|8�����U)U��!}�B�|m[���cq���z�$߈�G�WOF�>�LX`���� ���T떶6f�{�y��G3����sRXɀ�-p�mFNY��}�����Iw�{f�K��{a]f��g�P��L�Ň]Ǝ�����`�@�4=2�lb���>
�i�b~�Xp��NrQTҭlX�Of��`nE����Īw��8�it�f@\�,JS���c��M�
h��y�a@�<&ex�l�on��Y"o�|���w�%���0 @����� [l��ՠ���@w��75����1>��ņ!v`�K�*��/x�
fx\�-i���w{]c��DE�:����4sλ<�� 6�*��V>�s:|L�'���5�(q�.R�ު5���y{Ŭ�z��I_�%�WwX$�3�>[�&Tb,�Ց+��M��w��ŀY�8����W��"���vo*|����������Q�sl>⭒�ps���^��B��~'��_�R� w��݀B���Q�l�Z��A������]�_�{��\����cI����.+�a�{��GX���K��z���W�����WU�41\xul��p7Ԑ�H�*��M� �z��ė��vT[X�7�Q���bvg.��k�T?�%�ﹺn}t5���	�E9UB�4��Ko��zO����CM*f�6�tg���/f�ˉ�|�\6��5 �f����{Ó��w(��r�׶i��c�2��^�G��s�p-^K5�H.���[6�CI�&!+�����!�֜���V�\��nhb38�&R'��0�A<�2[�I���4C�c�I�+5��G�����*,��G`)��d�+��@��r�_>c��w�uS��A��&̉KDG�ȏ۟�R(E�X$O[N���t�=6S{-U��ޱ����]s��nL1�B�Oe�	�*�Zk�D^�,
�8�&�����`�Րg�c�t�O��l�k=[_���zh~vWR�����-v����F� =��[�T�g>� ��;����ұoP��Y>�1?�~�E�՛��Gʋ�r&�*OD�Gi��j�����o\��D}6�^�����}��d�w-�K�\�U#z��YZ �3:IC�����H��Ed��?�FY�^o�mݐ0L�dp(E�.x��z��|LC�O��p01���\�4Ɨ����kj�"{����ሖ�#La�`�k�)%�*�1�yāE�x�Tf(5����2��0���em�y~)|�(o@���W�(�N�M����5�1	F̫��D�iQ%���ˌQRQ`2.URg0�V��`ښr���f��m��K\}'����Z-�$0�hp�8�_r �}�N|&5dF��Ґ�k;#�ɑTDg�ނ�Y'�`�|D9A�f>�����®ճ����K�p���)��_m�B���7�	��
~������^-�{@_�l��Wa���b��"l_"�"*^��yb��}�����Q����r�a�qj&���w����ا���f����n*l'^̮�S܄	?���)�f������C�E�s��"�ofWJc��$($<�5[s/��K�{&�o#K*��@q���Ag��G��0��đo�1(���]�%*.yg�cu��2v9`)-��� v�dƝ�Y]�T�FS�'u��Z*1�?���ʕ�-2��:X��e�KX-W����k9v�Ư(�k�§^�)ǒˍ<�hT��#ɉp��֋L�q+?�e����I���Vႉ>!K~o�sFP�=1l��\�e�=�T�9G7����К�?�	TD��������?FqaYk�6kW6����~Bܾ�g�ɷZ
���$Ό���k��e������L&܂���T���?��T�y^�5���3�eZ�ғzD�;hf[������8�������ۿ�&�a2��o�p_>���_T�
9�~X܂ȳ�o��)ӷ2&�5~�ܽ�4�/T5�C5ỽ��)]�	�rSG�'Q����2t�{�}i�|s�8`��ΪdD㷥qe��Վ�x� c-�U~ݙ�*���������|Sy�n��.��+K�1��!�S�_[������������d��\��dBNy�gЫE�.%O��M }zP�G-���W��o���?F% k�7�,�����Z!��a���������:�6�n�ݲ��|�s��t�C�k�ybe�����8��ݢƘt��QVPeTO��:Y��	ϧ�(�\Ֆ7�$�O���^�O�K�ꋡn�S�*Wq����ѧ�/�тd�
e9���9�	�K�����]E:L�����K�v�~E�͕��LCN��c�GO~$P��ծ�����<�Qn��OY��+�d��rb߽���c��u���Ƕ�e�Tg� S*d���>dX��_�)�����Q�>�u����]O�UB:�����{07�ת�&e�a
�F���9ft_W�x`�FT�E��͹9X{�tL>o����Z��u�lk�:8;tI�-~���x�s�D��F�E�(�E�$�#�`p�y�^���OM3_���I���x�[�����b��&��)8����|�i��g$����
]ȅ ����_������ø�# ���r�l�~��t�m�/�.P�Eu�l-�xd�u��I�p���kA���?Qo�v0
>�9�D���Nj�}Ixz�C݆��Q���A�������p��aʖհ�?�:�x�)�`�g���n��^ Rca$��D
.�!(�
E��nL~�D�����O?{wo���_P�y'�e�1u�=�_��i����=j���%�wm��}�(��)�n�ޙ�G>��j���K��2ԛjX��+�Pb"=�E̽������
��t(X�W�#��v�W�Au�w;�x>|J�:���?�U�~�1��O��dxf:��8��/׮e���iu�O/U� h�w�U�Q�5?^l^�I�a�V�_ �{)�B r	��Վ�2Ay(o�J��񄂹�ñ�#6g��{��?�.]\
oD&�6�>��j���G�+�r�ߨ��(�(�f\�H��N:vӃ��m�2_������C%��t>w
�l@&s�X=QP�>��a�8xK� ��������Z�;�����ϋX�K���B2�x�9��_o���ܥ�=��4bO���.���VYS���dJ@tB+� Rt�,Yɶ�m`a��Nx��J�\`
�y'�T�ԵJ��z�g�nFk΋*�,X��W��� ��PdN����l%PJ�8嫳g߮.X�Ko9�YшsYdi��|��d��	���1ѩ|!Ő�t*O`��药+o��Y� ��։E�{�\Υ�qe]�����1,0�6E�h��P6�ެ�x0�)�m�Or%SV;E�6���[@sa�P\IrB�{^E�h�\U�_�-}�&��~�T�
���Yw������Y<eչp���o����I�#�n)�jt���6�����=j��#�b^q4�ڬ�oR�}��[�cU��]�dV�g��|f��h�v�+��l���f��D�A�Z�0mؗS��lyih,���e�d
3FJm;��$����G���x4x�C�Y,�~K��������알�U��/%�S&�i�l�P������D�h�K���2�����4��'t�}�ˀBQ�V��(@F�������Sw��e���./MTP=���F�i��������S�E�_�5;4o=���9���a<?���8	��}�,|�l���ޙ�
"Xv�x���FG;%��(>�(�&L�gRa9�"��!��G b��"�p�����'���͍�8��4Fy��c>t�إ��v�-�i__�_d���I.������R��S������������o]{��I_%-���gV�(ţ�����i� 
��'� �۸��1+����]�K�~,X�j*�`J��=�h��qQ��
&`�`�l;8X�v���,0���
�}�҂�Ť���=��.�:�bB�%�PZP�:�J�F�Fփ���}�%����]�vۋ$%�aw�����^�S�[� ��ǥ)0m]��0���
�P�eq�3y��Q�x	��ٌʅ�s޴G\<��~�����(X�+:]D%�F�PF1j�I�A�  Lm����~V7�nmk4��Qg����G��H��:p�!���&��9�_W�U��wQW��qQ���� ,�'^
:5����,��=�$5��Dh�wa����_I{X�����e!kYӿޠDX�����W� ^홊���o�x��D@�Bt�Jy�&�@G#�؝+_�M�b�Y%ؖ̚�'{+_���{^"��}�YV~DL��I��٣oEX�Qĥ�W&�����J%�䍑0�_|H�u�4�^���OCF�����4��5�������pH�H��[h���r�*(`uݍ
'����N���;5)�_���։K��b�H������y+��0x�L�F8\~ �@,릴�@S?\ҳ��5]�"c~�5#DWKZ��)�sI�����a�F�� kPY�|R�R�pԩ	��4�ѫ�`�ll�(�Z,�Z�㚣�ڛ�o������Mf?�C+~�Its�s�7j�অ��8�
=�uGu9B�ی�yc���A��E��OAt���L��΀s�´�����x�G�7��{�|kĬpϛt�١1Z�0��Z��]��n}3�yIg�.y53��o/�%B�v�4O�ŗ�����eHE�#�fNP>�L��<�L1u��L2QYU@�
�!��וxX�ޠ[��Rl]�������T/����(j��p������ʕMxMS�����c��G$�Z~g�Q\�Zv4?l�ك�
�L/�{��� r���u���5"�sn^�HLɞ�'Y�Z~ew�_�+�	�C6:1ϛ-n�;4���8��6%ħ�_^e��p4݂��h&9��e��Mt5aE6�Y��Ph~�����4Mq�}����@ 9҅��4_�󀥺�g�.�^؏ʳ}����l� d�y;������`��}���
��
a�A0/p�,fd���f�g�s_\��f�b����E>š���l��'�ń|&d�q���g�-̊Ս~ou�vC�SU+I��)<"T+���[�Dd����6�WS���&��vN�.�����y"�x�7J��V����]�RC�3�E�D�$d�����>��w���<'�\�֓��m�����ɰ�@ֹeZ{D{x��].cO(eG�L�Q�M;d�[|��FJ�<�������E����2H��C���c4n���E��Ja�M��j��h��1@@��(��9tU�s��?>&�3s��3r�tCw�����o!8����^>^p+���B�<�?�J�u#zc�*h2�!E���7#\GR��XDPC�9�Z�Ť��?Yf*���K 3�Z/=�%������q�"<�����󫁢�a� �f|���O�$�]�-/�����sЛs�rQ�k%E�l�?
�dZ�1�1~/X�e-����%���%c��D+IK3vAA��0�d�?�õr�����SZS��a�:���7�'i�24�JuF*�dw3_3⠥�֫������G+z����z����!?���xt�0W1<��Dc��{U�^��\�?���E
J! i�|����ɶr�>%�ɖ'PM,b�>1h�v��4����)��_�Q��$�d�M@��W�'�<[�H?��{3Ҥ����;���-��>�y���ƙ�J����Ey���������ti���=::=�	=+{:��-Z�r�Y$�b{ ����i�zT�h$>�V���{�����2�M�^6p��$�2��8�7�W�B��S��eA���G�; 4f�>!�m�e[�^��_����JG,�5G�yU����@'@�f0��V���=����*y-�AW�X��U��q���K*���$"��� ��$ս/�P���#j���͝F7�	S��/��5g���7����8���k:�!��nD ��z8��E�D��<2�<����)D�L �izP�Ͷ�l��hw�� ��+���#��>N�~5 dĔr���m�L�r�J�.��MPZxyC���F7�>���(�(�G�~�ŋ��4Cy���ۿ�8�v9��
 ,�,�DbfM:4���^���K��3L�j�!�� �%�����բ��$��^�Q����>����M����A�ǥ{޾Oe��{^ �+��N9w�6��c{U�*Ė.��~�`���\d����w�Q���t_�Pi���gA?Ѐ��)�'�4��Q��P.^������vl��N�GvM����,^��)�\�m��_��6�ߜ;$o _�1�o|n�@X]�  w�H��EU!8��ܺv�
��?�[�e�P>�+[&a�E3CQ0��lta�g,
Ȫ����j݇��;��%Y[��s�}�9����J�F5�lcB����:����_�ֆ�΀�b#���.�:����x��#���Ő}�g��/�SQBs��<'?D`���L���gӃ��:I�����I�?:���u7�f��
���? �_R�0�ͩ�Ԡ���+�*� ��2�=�LG�
�U&`P�9&������h�fٝ�K�«>ߓ�ch���ƭ�f�O���I2Ϥa�aͳ%سj�̹��Ƹ��\��=��4�e�������VF�P&h�>z���>�C��^��7�����[������ZR�.��!-��K���Rp\��QH3n��Q�-�WNQ��fWqKg�����3J�)��`���������E>$���Y������ ���>�̩x3,���-g�;��>'��)CȝnK�n_�׋\z`��]�}��J�5H���QM]@�[?|�TL�}���8�,$��˜KuҦ� ���BT����έ)U��a�?�G������	_���d���4�����f��.���o`U=�l��OF#Jl��n����3���i��|P��@�k�]�Ş�w�OmU��{�C��ną����B�d�m��r��'3l�uY�λi|g�M��-I�9W�����2�4�'�Ƶk[��b:"l�1�A��Z&&�}G2s�*�ʡL�0�L�����o�_y\�%�}����:���X�2����\�f���2��t-��8Or�[����dL�0ԟe=�3�C!b�=zS!�
�� ��cG�8=��]�"�*�����{l���t|r�N)�D곃^�+ۂDVh�|�t��I%a�q$��{�n���=ٜ�>��+�>�q�@k׸�)�:{�R�[]�[��ݘ�z�a2�o�������K��U�'Uuu�G�̇ Q@'��]�g�do�)O�"���ӯd\����.Q�:H�F�3�|��F���.�]ݲL�B�!��Q�z�m�2 �{kOI_��+���b����KuN�c�7������Qs���f�� ��U�@0�n�KCA�OҞ�)	����9��KoMTRK]��-g7��F$WH/K�c^�>-Z�KA�MY*~l aP�����m���;Ӫ��"1
v����pV�X�jO�zs(^�����r.�t<�����f���i��������2�= �T�ϑXm���-(=�[����H�r��?kI";u���`���.֒�[f�����8h������"Ϝ���Y;��\�luvM�g@ۺ^�q�u��pk_��G5�AH�C�Yk�l�|�8��~��G62䘉��i�K���Ԉ�!�)���ǐ{�P�L��,C�1�v�_���ɋ�_�u�(�9�.:�<�ض���g̞����g���z��x�~�o��S��*U�Ǣ�3���6�`����˴�!�!�����7$R��}%^��g��&_m�[@�����8!L��� �u���c��`�(v���!=%��k�"�q!=l��4݋�T�~��K�SeV�` ���*�yQ��[q�T��	ʦ�ay��z��d���J�J���A�x&�Q��ЦN0]�!�69�<!yL��ڹ�+qoO�\��Q��hz���p*>	8Xd�$�i7�Q��ȼ!�,r,�� H���'ωZH�%��a��9s��7�ʜ��33����ĎV,��>����I����(��i�������5:G:N�$}�[�����Ծ:��c>f3��5/��SK
�(BP ��� ���q���>@×��N�2��ͭ�0̾�֣�����檾7���p�W"�O��Aқ�-@��O#�>��x�#��q}�r ����1��	�v�?��>e䢁���v����"��~��t�{őo�M����=?���)s�E�tH�V|jWP�1�������,���P��4[�@n�Q�+��T��}'�Ik#>��0�T8{nr��$�X�ׂ/µހ-8����Q��P���J�f�.�62s���S�`= �hxҨ9��a{��Z2
9\�li^ٙ������m�\/G�D,����mDf�YxV3�i\�fVY�\�Z.W@a��}sQU5+��A[�㡢�G3lŢ�� ����NU�f6��n�CI���V�tؙ�m�'��bv�5T@|�!4F�d����x��k>��+��<_���n
��iS�S�6���?�˳���ưع+��X���x���O5�Sx��!�1֞�����A�ҨcJ88�  ���q���]�J��%C.�~�BGn�f=x,�\�����&Qc���[�����Hc�v�&2|A»�|Y�� ��$�,A�;Q��Q?۸#���t���4}Ȩ�}���(Og<*"�y��ɦ{��B���a���������#g�T��g��&��sqU�C�4���/�?���J���(Z�a�q�־�G��������u� �"�E &����!��/�����c�)�<&�Y�W!W8�fj�*t,��73��܂l�q]׸����u�2�
u����F�2;6#��X�T�>:e�ho4fN��#0���h��/�*;Ip�Z��\U%z	w��M��I����Z�Sޛq�I�^ǋ�>���{�-��D�T�=!4�>��]p� �o�x�'�m_C���+���%ÞˢZ�aZ��3a�!�S�� A�y�nCzN0�+���i�&�JR�%���8,��?��D�)J�La�2Fk�#~?���h~q*�ΚW�%���U,e�}��Q�p�p$�+�S}�
ys����ptX�5~ �=�mfS 2�D�_N^��T��}�bmC���n�2���|� w�	����X�!6\H�����KL�Z���)�ȁ��d�O!�-���NP1�E$�T���9�v4�І�3��,���)�����q��&��k�,��@1d]���nS���9Qm ��#�қA+��6�6�E�Y�R]�$s8*�¥�軖l��+�3����K}2Q?"S!��ٴ��'�<ȥc��[RK���@��9���%7H�O��ت��`�D�� ��]�k������ͪX<���|�� �[nn�¡�qLq~�Z�qr{�,�L��f���qM��ILk!;;�YR�C ��?y�&��a31�lg���~?���i��1��gUq�u7��fg��	���a�y����Ge9��D��W���U8L0u�9����A.=R�#;}��Bëi�1G��{���.��n��ma2�Ww�C薧}�D���7_]��f���0c�>��X�䧪��?��R֌QL��+��v����m�f��6�Fo��.k��d ���ǆ[YUyV���[�v��*�	�3E��#{ར@��X����<���ɇ���8%��%��b1�YTY�%���u��r#�['}�lޡ�c��;�A�ߠx���jm|��
<�$�*5ϐRޅq^ ���G��j~f��Lq�����J4ރ�����W1���3�MM7!��su�}wYB�*7��kڸ�-껗������JY��9�q���
���C��BL���0<ڊU�p
��y��9)�ɟ���x���#�i��P�m�Ϯe��7%��{KN;q�(r�;�L-�SGB=0�}�_�u��9����?F�O��z���c-M����X��য��ۆ0�o���x[���!3�mV�Ӹc�-]:'�D�6��SF)��;�Y�z�r�O+���0ڻp������1ލ�R���@xxُ����!�?d��ϟi��	� (��X�\(�`��r
A}t�~I��qY�s���s�M��HD���$��!I��2dHUMoh��R���I��ߌ���y�!Y����?8�:%>�<�D[*5��oG���.h
F˞�i�U^��s�f�\���|��#���!Kk_e��������#Ԋ�e����=�����h��K�O1&.Q"���=`�8#�a.j�|T���a��:�����P��;K-؈��FD�e*L��<y⾎U�|���:���\k&�C���4T�r ����s8�/�/��Ha6��j]��޿�pKъ�BHإ�$��^ᣯ�6�,:�d�V8_�7 Ix��Z<s����e\�m�QL0��=P�E\C����M�N�j�5�6^e�Wl	��d�mGMT ���������?�(��;7
v��r:y�4;�3I��)ِ�8jh0v� �@?��@�ڧ��ۼKb}R#�3���[�2�vSBh��;��b�ZEJ� Ӂf7�cl�{_juJm�My������!�����)�Z'3�H�~�j���I�V��\�jC\�EH-��b�Z�b���C��ϝ�tG��z�`5��"h�(�����xTq�;�z�2��� ��Rv+���¢���7��d�&:�����[!˹b����7\%A���?�X�u��T صO���	/9���m�h�Z�^�z��2Y5��P����(��糢���&];U�ST�'0+��N�of�Tۉ���<>W��ݸ�!,�(G��FfF���O��J�?�o�z��h�Z+���?������ي�6��s�x��]{{H�	��aMK�f�A0���U8ā�h�>���xz���+�3�1��l�5���?O�7�*M~YPhf9�2�(zW��i�	�b���a!]���[:��.��n4?�H���dIM�f�0?���M�'�qazvk�����d}*C	9N�w��j� 3��GW���ʲ�f�����if�5���-����F����	"�}��O>�<=mR����_�O�v�7yc�P@u4ȟ#xLF���e���qnpݍ�T_�1b>U$/��c���:����g%�����h��ɻ�!�*>���;6�#�Y&B�&��MP6�r�52��0L[�,�q�
7mq�o;��q߱%��
	r��q����@z����<6/\3�I��+�SHuT��/���G��&E%.�l[
��ؐ��������Éd�! ��$�)5C��z!F��Iq�I��w�Ȟ�!)�i�s&L�i(�E����Sغ��pX��+woT�s*\��6�0�j��X#�,{7�Է����}A��}i�����M��D�-�q��`0���g��sK��Z\y,�����a��\�#�6���vu���aX�����'xj�wO��%�n���YpU��:哠��[n�N��LQD��^�E]���4��5O�yd�.\�5%A���*A�99���A�P������#Y���\�B��G������?z�tt~�d�ӆ��VT�-fH�)~$$ai覩@�7����х� Yz5\��%l?U�&_ܵ�����O�5��6!���*m�o�E�SuH���S�sCq"K�Z}q���%���}��UÛ��2�;BEGe��\��2;E��_۲]�'�Cx`����qK�tV'���Xb���k��S�{�g�~�)4`�F��(4L�Y���Κ�#�8z0n($FNF�uc���Us l��[cSإ�����������ZO`E/��eceʍ��I�z�獘n߬hVW�'��b6��qe^�pJ����i]&zI�kF(h�8�8�M�߼X���5�����lX��݀�}��O�+j��@z��R_p!��M��9�;F�y��6V.�L����������d��W���3g�q �6x�� ·]κxp�	<&��W#Pf���HJ���v��!���(�eKԼU�vm�Q�p�&������{���=a��o}/�t`���±�"������q�,����ު�H] Q6�2#2d�����"A�����Cз�|���4W[��
<�4q��(�趋Qm�vVw���R��B���@9�>(�&+Y��jt���r"t獯��E���0���<6�:�?�9��ظ�&y������m���r�b�G�^?�U�bci��~��׫�D�Q�����y���
I��%�21��?�
p�Lhs֜��}�uوY������42��a�[Z�������vP�(���t�^C�}1�JI2�ɱ������ ��R?�^Td�΃���@����]�w&�歩�ļL���_��,��-X���2���3�i�;�PR$P�D2{�;߀���ʲj�`kae�$��#�C;�X@��TU؞�E�U���v�h�3���R��A_l�l�	��!�S�l�:��������#I�@�?`�\'<��7B� 絩US�Re������D����J���6�2'��_�Ő��bc���ˏgy�Cn4+����g�~-����D@Aޤ
��8��T>���=6X����c(�^�}��}�9�]Zy�x��hEkK�L>T����J���(��I���ƍny"~�7- �rZP@�|���1ɠ��r��rM�o�ʜ�	/��M��_T���Hɺ�e�ߙ[�y2�V�٪0a,ݪ,��[~�*y���lWm�+��p�ɚ�`�ed������4L���e��a3%��� ��Z�˄P_�?1��(N�Q*�GU���L�B��������<�������9�0)f5sP��"|�kT�(M�o�`���صAB>Ϥ+:h^�����<����b��Q�9�饘�*����7��
�MV��I⢱�%�Qa�]n0��i����w�S	����ֽ�$�F�c��d�"c�ID����b(��	�~��{5v��)�ti�7����26��/i
`s��<��UD;�^Mx��:��|�W���)g�~���VKP97lɍ3� �'_���{����\�=�c<��z{x��q3g{^&:�f��(�D_�ot`-^��d��D�E�H:}i�h$"mG��K�9aw�$-h��<;���n�]�$�g��]7l�L��U���,�������ޚ�؅�/���a(K:v-1I�h�:�����j�uS����ȭqm�7��������@b�w���qEդ����\̻=ix�Ε�~&9�N�p��bR��@�;íU>';��3����Bc��#�áI��Ѵ�8A��.7�d
�ެ���_�)��㪂�|�#��
*\�#��l �v����r4&h��>C3�h��B�2�(B���jFBE��u��o=��6� �S�
�%�PɄ�S�I��H�m������Ʈ�섲$�a���c9��?K���w
�I$C5Dj�¸�gS+��\��a��Y-���d1iPiS�_�;�����k9([0�73�1�Pc����ӪU�k�����I�[5�D�8i������#~ Ȓ�-��LU,���(��o%(�f��Ľ����I�*C|Kč�x5�ށ>�;R�ݤ�T�D��>��{��H����8;�׃�p�?T_�־U�(�>�ܒ���hE>W����#���1��RF�.wz���/����~��0�Լz�_ ����ώqkiz̀=���y2:u�ʔ H��DT4�N���4�
�@��w�2M �b<�k�����?h��� �M�Z���a(E���c� "M��7�%8�p���3�͠+�?8���l�`����nU͙_��|ax����i�]5��+Z���ՆM�P��-s|�7�}�:�(�1����a9X<Z��� L4�c�e�/��f�ؓ9�+���/�[�B]>z��J�B��k7�1j��_+����*�F<�d��<
�yc֥�R��
e�Z���G,�hXba@{�%��M�w�Ɯ��Y��f�n[��W��kn�}N�
�k��ާ-��<c��k<�	�-F٘@�Qg6[�V�=?����u+��L˵�Q�G5@���8FauZJ��w�_"9i�N�f4 vڹ��>�k�tS5h�F�Z��%C\C��q5��4�
�U�+<LN�����ZD�����oߴ�0�զ�T�����<T8F�_L��_ ߚ�?F��Ў��$IU�8�HɒF����3���qNL���b�"1&����N|��;�I����{H�N������ڈ�a���=Z��Ugq
��r��}\hE^D�u4��Ξ�i���f�}��_BA��a��T�9l &=�s`���f��
��� ��e�����FH�p{'G�텼�vJ�)�,F!��a����A��,���sr�܊�\�y�����=tÇ/�٫OJ"�����N% �$a!�{�/�g�����fo��Z�Om?��Kp�&kF�N�WDW�6��_�h1�>T¤�Z�p��xul����L�?ѷ�7+�k���vm����I�B4�Z���Ϯfj��A�=�**�r5j�$������d`����u����(��CC	��;���J��VDu���7=~�`�����eI����_S&�+U'��U�ж��Xdy�M�d��|��4�������8���@ KJ8��4V[�� s��q1���O�S83�uUiB�h�1��{��Zb����W��B���dO^#{\�y�i��?d2��`5�	�_p"�T��v�]pd}�=���H�pq$��"6�|X��dD��C����y�(c��ꊖ�&L�mۧ@  �b����ji�Q>,�.�s�l��!-M�n�~"_�is�R�@�gW��SL���.��薴���\(w���C�
��0��9�3x���c�h	N�O�pS�g���/2�&�?��ˢ�����v�7ڥ��7Nj\3�kw�kb�fH�;�m\I Q�%Ŀ���]_�	���Y�q�w���K(`K*�)'�}�W+��g67�)�ή�	~+�8���@˲`;D)$�'vCrE�O;���>�g�0	�[�� [��^?]�`��w�Zs�	N$�.�+<m1$��H��Ov��Y�X{(�5�!�	3�7���#�2��1��-�Sq��H�� )5�hN|��8�Z~!zJ�����O�P|Ә& *�X��`�m?�4�c��҆<��B�v[765 �U�G���Iq�@P���b�9wCK�O��#\g��*�X���������>���7�cR jBb�H�~˾�����_��|� x��m�᮲��F���z�9������J/5cdD0�%�xW��z\$�|Y�>�ϣdn�#�tP-�ÿ�ȩ�q%��
Kݗx�p�_�ְ��z�qE��Z��:<�N���Jc�t���)���	2�I�n��iȦ,a?j�f�iBZ�.��!2� =.P��x2%"ڑ�|޴�rL�Í�RN��=a�?B ��;��:�oh���He����-}#fZʨ������3��a�e�l0Or*qD~4t/�� kA�8U(ۃ�g�C���{���8�ߑ)n5�8N��� y�~9K��N;�&���nE[2Mӑ���s�R|�O �8I�"Z��-�<{]~��	������4$����I�ޜf�{��x����c;�o|�U{�_�#B��u�x�	�$pWϨ%&���P�(��SM5�C)�����1/ 2p.QW��ry@�!nV�NC����(O��NCb�2�	6�h��;���x�X��ȫ���F��N ut�p>>/l�lGT^�.b����d22��}h����ݓ��R��=e&�ۦ*B�d�s�4R��ݲ!������(�e���d�=m� !&4[A���Kh��m�0�ƨ�^�l�**	G�,b��5:��Ⓢ`�5�B?Z����H�'JO����q�����.�0l�^k��&W!�����s��)CT�ǂL�|P��C��꿊�R�[8Kd<^��s��ǟ�9c�?�FL)�J�toA0�U����g�Ոw�ܛ�y8�}ҟ����-�u�0���$�����(�4����R�>����{&�krSʚ��,i�������W�=An5�Z���z붶fGg�14��i��+�v����g�jKk���0s_��#�HI>d �W|�T_vxI�/�FDND� �v,Pe��vȆ4�5��A�R��fs�d<���i��dȲ�cY8����7��
c��@F�#ʬ��M	Q��lӛgI'�{�u���T��u����4���YP�^J��,���R�z
�u�A��\�ͧ{9uC��e�A�v4�����W{�}n�� �;s�V�����(�i3�^��2�*~xD���0�5�k�sЭ���#��7N7)m�g�k���5r�o���Y~����6����Um�֡������K��ܫ�} �����]6��(��A���pdG�<=��飞'!��:,d��*6-���VlSE>I�Խ���3h�L��M	Z>+��t�K�x*w���[k��Fҙ��80d����V��n�p�V8�6o��'ĜHDB:�SS�v�@WF���$��[9
?��D,�A;�m��q?1Duq�'Q��'���xކb%7q�{��n��_
�~l��qI�Z;���M�f@�����}h/�f˔�g�ig&�IFض�����;���2�*LW[:nu���oV�,���=����'�r� �$�oӈ�6!� �e����N3���?�8�E�t�������a�9^���H^�q2�|?�(�ǬH4@5��!�;V7�L����C�gˣ�M�.X�T�����r������Ga�o-^�1`_׿xk��wBkb�sU�U�lV���*�e�^��ρ�q�,���4��%׊���f��k���j)j �J����6�3��X�~fy�����;kS�7�����S��H�r$�8�����a��st�|6�#T��d2�H~����8�oJU��nڈL�{�I־_^����,�F��=�8-��9�ρS\T��2w��4F�&
�4-�FϪ���`�5c;,�dutd��5#8�^��`��[��� B�&�'�v;U�u����U�������*��<�ծqO|��WǇ��7<|��*?�!c�����U9�E����F �I����qu
,��J+(,���+v��(`6���q�њ�8d�0�ke�����$�¹MW�����T�%���(^��J������12�zr��e�+�فX�V�vz������Xs%8 G�}�Qw��I<6�\�,�m����^N�_�Em��}���[��օ_��a��|����8P+VW�Uѐ��u��z�}�i�y�2D�2ڧ��X�cpd�Up�|�)�b�ΏR+X��i�k��d�&Ml�6u�v�Q	7��������K���
�ˇ����V��e���U~B����� �W�G!�Rr�I~U�U[�d�U��r���
�u�G�y�R*�m��W�6��SD�ݏ�/�>g
1���X�`>��G
�N�`��a�t{�Q��5[�O�6B�Y�h����)7R,_\�ɟpH���/��B�]�T�&w�w?��ަZ7�MI�����Ժ����b~s�5\qI4�
௮����hb�x$K�ʞQ��Lk8�#\�dW�9�����t�I�G,0�H�%uS)�7�2� 
\������)�lא���R|��&���s>t��Ue�ᾰ��ґ��{��ϩ�1�3�Ƈ���Z��G�X��?*b#��:U�B�����8���o�����\�ҢPܖ�QKYE@�~X�o�?��KFE�T�K��}����WA��ko�k�O�<���qU.�G��"���A�]�O�2:��-��@'������S�r���G�VG`��M�Dj_c��ZƔ�w�Ԟ#�����F���"�����Z�>cJek����Z�v�'��BȌ���f�Y�{�J�v<�|nf8/����w;)�&�?�N>�\�t���G)��Bƌ�4\Qs,G��Ī\�g��0�Y�
*���V���=�����8�_����	�ޥ.7l�_"��h��@#` 叇Mg�����x^��>�u����6�X�^J���1]w���X�W�J��9��o��)�a��#vz叩0��3���%��H�����ڷ.N���=�y�'].�b�]�9��+�y���P�*��<��9r*0�J"�I�������h$��h�Q���ʹ����Kg[b��4�P�L��uխx\�qK���R�,�po�^ ���4�h����.�]ȝ�d'�@rJ��V6mx���;�=�)B�(�ݹ�L���A6jz�O�'$���*��E ��$��K$�5�J���)�?J�T�iR�f! �>a�+w5�"\iǬ�,�������
�$L�Z#�q����=	���U�@�w�p�X�	lPjH�S&^����k'�,���j4�w�-,�1����c� /�e�ds�d{r6�,�a%r�bW�9Tt�7�Y�)�]�r(D�\��gH�r��̍�i�W��	-��E������-�Q��ِ\@@����Op#��5Ռv4��a����2*��0�p\��OXs��a2����R��o�poT
�m=�A�Fe�%��3`ԣ�ӇW�����V'W[F�-焑�o�+ZR�rWPH�Ƒ�aa�F�z��{<���6�[�l��[�cٛ��o=:W�U����zF����4����W��ɟ~�36�c��^���Ml��e��h�"hI!���,v��.Q��"'�]��b��p��{��4�Q���ڟ���F@Ө�=�e%F�u#k����X���4ȅy��)��KX�,�Y�WC��<h�H��Q省ɜ��t�6��MvA��KiaPn�7�'D)h,�����V�@�LIW���`E�H�����jD�+_lkS�#�h����5-:-�7X�H��H��!QI��KeY�y���7$�O2�A�w��gzϯ�"��t6��1d�18E󸂭Q��}b*�5�E��+�&c���G,���.7*SIp�/�����X��mږ G	�\�"���G��c�$��ԗ�J&]LH��B��.b!�7�.�X��܋~�F=���Ӫ)Z����ք%' �OH\�3���J�K�0c��CV�W�k��I��@�MV��px���D>6��F2��l~]$�h�
&>��^N��2�@��jƭ�D����Zk�)���o��|��c����e�����5Qf ���<�y<ʯa����S�]�d��G�]&�d���r�T(=ρEV�0-J}@k�m�Z0ca�O��oRX��籅�d��+=P��� ��[�I��t�@�܃>������9{�;�?�Z(:�=���P��o�Q�o��o<��8�*�Q
c+1n��BR��!,Y���S�:_
���S�:�dE{*:B�:���9u%T8K��RUNK���O�v��LIq�r�fw^������o��X����x���N}�䉼�y2��g�l3<��w�+���;}����A�x'J
h�W�@�+�]gȤ�q��RC�$�<{����5���.	U��9"��}��{]^pDl�?��e�u�܆MN�j�:G�?���F�sA;*��)¨� v�C �6mıV��MS4�}���g�o&�^?+!�%�g�1�=��[ݏ(��@w��.*��,��_�/.'�7w♔6�1��T������\��Ъ��Y�}����>0F�d���s�=�L�Hh)��@T���Yh���>V^L�����`�t.���[����[ĭ!���D�jv���8'�n��#շ4=�>���v���霥��ai�bi�`�������ޜ)��D���f��byl���8��[�ǂi^��gU ���#����{]�[����%��v&��jm��t=�V|�ʧ�9U�Q�#�v�!x|��:c��N|�=kɳR
W1X(� �r�:'�+):��+���qx��r&�5c?�ʶP�~Ϸ�f� �Q��^R,Gv����߆�V�X8�!����5琥~s��}a~lbMV�Mx!0p�@׸"�	�kzv�+�?�́q;�s�9X�SGc��� 3�ŶK��F>bv
"*�����yjԸ1�օ}d5��ۭaDQ4u]^;�i����#7N!K�����1g���4M%���!["yhx���7�81%���_���X ��	�0E�Q@�r�m�.���FA[y7k�����"�1fhl14�{�GZ8��E��6uN��	7,��j������A����=8Y��v��]�{*�b$4�?���m�a���ږk5y�<��>> ���d>�>��'��
PG��v����#��M��Q�XL�iS'bY
��	�2r�s����"
�-,��z�q|I�L֙��83�\�*;5���n�*���w���ڊ�i�~��~���Mmz��F��Fѐљ�����G,����(���h��(�����H 3�߳b3]����4W��Mg��Iˊ$��d��8���r�w�O�pB�x��)�³c��$�c��Q!���$a�}MN�ԩ9��_��1"&"���,�Xl��ΈC�Fq�F:�잃U�u�k��@*�b��Y�@*�8��Ky���,'��Dh��{�p�=��g�v%�o�̳��9��Px��`�_47��)���j���2�F�a��o������нr�Gօ��a��.�*0=��E$G�r��ė?�9���;�B��|��Tx^�ú���?w�4!\1f��׵�����E�/�B�?$�=�ˣƶ�"�ų��^�R�Ô�Ԗ�ԯK�r}�`@��.搘��UE?!�Ql;!3������C�����P���<����,��6�D�cө�e��z��C��a1�M�h��$������{��Dk��z�Q��`�`����=�T�b���tN�dm�й]~Rф��f�zx1�T�`���J͡b��"��!y-�<�aS�
Qtъv8U�O~"*=I�.����`g�nX����p��$Zz}��ּ������p2�:����P,J���r���8�@ὦt%�y�<�O�v����Q��k�K ��!���޼MӂGKf� CLH�4�,=;�ǚ�ٯ�v��!~��)P� �.6?���A0kS��������\k�?�IB�0G��+�����:��5�S���RT����+�aJ%���K��	k�TS(֣gp;����P>�#�Z��Tb�1����O�N�e�3�F���8����o�{P)�P��FK����AvFo��+P������-p\pC9Mg��%����u��n$�{¸W7��������ZU��5aG�?h�%�b�j9�S ����G��x��{n&�@q�"��-uF�$QF���MR����ڇ�F�B�2M�L�]J��h8�e�ce�]�	�����TN�$�f�0���>��}��U%ݖ!��.x�ZD�SX����"�!^2
�NG�4��5�A4q� تuz#G�
㰓]�|,��o�W� C���-Lr���&���<�9T���ַ�w�uU,����%�*�g���+��q-Q���/2�W��v ��[!������8��l�қ ���h�!3�5�:����Y!��zn��T=��_�v�l�a{5�q�M�	�ԁ�N�[5S%���@N��J���@ ���˸��N�a��� �7۷�i]�B���ߡ#wH�L1�{5|2m���ݝ��sqc����Kp�cp�"�x~`����^!�1�.V�����9
B�w�~{ˇ������VZ$gu�����<�9*�SQv�"�`���%}�"M���:������z���3��0Ț)�H�cnm��L�9���	#�h�m�x���ma�Kk��l���"��E�ڝ��i���Ջ>�Oݸ��7%$�4�/0E�_~%�Q���j-�"3�/�e�ע�1�ȃ���ݡ�@���ڝK������V �u�JA��=���vZ�d�:�؄;ld�0L-#*�=x-
m�85nl���cO� �x���F��)�^�I�tM|�!��a=��`~�u�W�$ǆ�����3JӀ���wPl��&���j�\�� P39w��Y����'�t��5ۀcw��Ma��)U��l��u�9���D�<G���Ԉ>����&�M2�VÑ(��C�]3
�����7�Z*�F�mi[>u����1�w�l�w�/�!����S�D�:��R��!��De�NQl7�b� ���Ⱦ�<gz�l8?��J��i������.z͙��S��2'5��18��P���gd����]vh\�2�@�ky�_%.X�$\3/W�Jc_�X�$�����5 ��,�& ��@+����D�ȑ��8Z��m��`V�
��Aw��H^�b`��z:�w���*����d"��T�=�N$��T\�Æ�(t9
�P��o;U�*��b���zذ�~H���`�F��9c�އ�w`A��3���YuF�EQ���h=kC�g?������ɢ��"+0(�c�.I�?��C@|��f�X�����ߙʸ���"&���{�6���8�P��yT���+�}��"�{���rѨ��,���3�E3��OٳߡN%}�ŠsL!����̐�r������L�d}�sFjԯ,η{��M�"��	j�Y�<P	V�z�9�Q�B�� u��D�d�1��.���Į8c�h�h���LU��V�w�'�����"?�?e��K�_�f�j�0gIGo�7�<�ZB��Gq����vE����=�L���W�bH���C[���C�W�i����Ŧߥ@o�����ܛ��8�������Qe���w�'��p���%Feq'Zj���v}��"�D���ߵd�܊�V��=>B��O�^$7P��]����e��9�˯�j��U�d7��� �V�#��0��������(�m���x�q����@?}����	7�@������\1&�j��9bl<Q1L�^<���_�M�� �#�O��i�ѷ��Y�ș	T"�KƯH�ն@f�SZx�a���}ܔ���B6�ުq�	��"�$���'��Q�`{�F�y��{���'�V��Hw��,���(��x}�}	ۆ�h7� �p�g��Z����0Wu ���J� Sߘ	����.u;���8��)���pX'������0�7���v�0���e��u4k��9.*[
��b���v���g�n=�dG+'�g��0�~:��N:����@@����lsV�\+{�S�
� ?1H�*� ޣI�x/��bX�t>GC?���e��7�G�<�/�^!G	���7f~'��_%@�(�����;U���G�NIP5�Њ�?�t ��S�����R��|ՐT��J�� ����p%ε��@ݏ�8r@�U�~���D^8iC�c9 � tjvn�����ƭC��E���Q5�H���+�y�ƨ,��6���	W2�f�z��X.�o��!���C40���_�z���5jXC�?��Qt���5��L-HgL|�WF�ˊ��E4�M���m������@�Q0=���־9�8$m���P�%�'���\��r��1�C԰��K�;/;�I�ً`=�I�Kjp�W)C�p\�X��6`�}_5�o�^sz"U�A�
�Mr��x.��uW�6�U�Þ f3�w�l���QO�p)����m\r�z��/�%���>�Ds	�]�"ߩ\ӟ �;��~ҟ�p��i���Q��ط�V��VY��3{���U+#'q*�506p� _��fħ��V|�W��S��QL�"#1m��%O�m#��_����jN�T��e �[�) ^�-�i�79��=��7�T��� 7[�kt���cnFpv��B�������#W�R�cʽ��uȻb��6���}ˑ��<��Ho2/1�B���1����Pl5[	zsR7�R���S{Z�s��!����DbG�y�f��|��;C7�J�t�^�����){����2N���F�	���ӹy�7Q��V:J�thp5�*��HN��"c���kƀ�>�b���W��~�U���+�ALS@y��5�x?fރ���:�_�����^>n6&��g��R��������KMr@�B�-���j���p-�՚��|�����Rss!�VWP_6F# ���[�5�	K��Lt^�N	!m�^���жI5e(�=G��ʇ1v!R�g^�ַ]� ��@uߪ[���Y	m�y�q�_(�/��E�y�U\j�"tJ�����m!����n�z��i���yQ����R��@рx�)
��	=���-�^����3�»e�19��D��5_�/W�]����)�!L��PH���%�(~W
%�+��s����.�M���b�2Z�EqN��$����섙�U�[B��<R�f2%w3q���!��]���f�5o�w��Uve�����PG0xNteڟ�2U�F�l�RV� ��Y��vrT�&ߺ��Xj��YH���(Q����L!����d1=����d�ȳ��*��Wo�2jXdy<�˶���hW�x�/E��ĽPo襨U�8[ܽҍ�V��֒�gn�#���HYPeW��٫�"1�B����)۳�0Mmm���x7B'�9����G�+%t�:m�ڻ��^����v�}$��G���aO�Ҫ̓)���?~�Җ��W��~Mwr�fE��U�X��>`�1��⊰W��NN��n�r!�;et�>���)5}z��ٷ���n�ʎZ�=����~�l�h��y}�UFz�H��|-H��!�h�t�W�����GO����
��Zbŉ,x$���Ժg,������%�a�;���?����:?C�P�i7(j�c'|��D%��g�6/ٚ+��Y�{^0d�Ϋ��Vd�X�~�\I=i$�:��&˒�ƸG��lGwNx RԠB�7M+f�1��Anj�cOт�-� �$f(*(�h���8%#���ر�W�$Ϣ4�T�j!VsQ��1g{F)·�e�8�\��3;,��p�L!�ZF���d�eʺ�,��f��@�s�3�vSّ���2���ZЙ6D]�r�%��I- ��� Q����`|ѣ�p����6���|b (ĂKZQ�M�;ƩjsHy��@����Y̼m
:��|F%,~�}Rd����������6�F�]��ە�2��W�m`�'Z1�[�^NovSr�;#mE�< j�n+��ߏ�Aڶ&���{���_ d��D��]�?�R�T0��$\�������*�fb��}�MjD��
�4�	di���wl~u?�#�Q��p�/=�gnP�ȫ�����VZ��W]���wFnq�Y�1���+-{1���"^7`�~��dd�D���hg��|s�R�p��H��@� ��'���Pzi8nj.Df��/���A�|seX�!�4�����O�V�yu3����Ŕ���"�M��A�L\����/����Љ�>��Ȩ-Sm�k�~�.�����oǟ�F1�/2%Q�1��G,��Zᩆz�c��5x�����2��R������=Yҧi����]��E��)P)�z"X�dŤ�omm�^���G~g�'�=�pM��7[D�z�4��{_�����s��}�*P:��=C����Is,�lX��ﶻ�02��l�!�|�/:��[�B��I[�A���Z�P��CQ�|/l����O*���k���=�VݹU���Q�6A�{T�����7 �7}^��ɭ������=��g �?�����ֻ�U��wo$���d�9���]4�����g�ƍ�~
��q�
2s�rv9 ��^j�T-�5�=n���v�X�L���� c|����L���B�J��kޢDE��F&H[���Y#<)Vu1��q��6���J����ʦ�H��䜯�D��[	���� ��a�g��.urjgu�5��5~TPX{�|7��������'��5��+m�Ø����zי|�3ӌ��
Xh9�~�{)���ͦmb{�1{D6 �fM��%i]��~+� ���ЂsjEmx����iF�y5��l4�=q�r���3r�K���f�15�UP�Ʀ�@��뻨�!�8��E,
�&6�:m���O�^�PlSߗT/�vtQ:�R_�4�W������=��A��NeI��6�E�?ښ������{1*f_]A�h���VK%��fJ���➞o���]P���Km�#�c���kk���O8��B���=>XQW���(�*΢�]X�Ybs V���l���I቟�[V=%9ҟ�����a�v�$�{�TU��5�a��q�'��Y�5����z�_6�9�MӏZ&�Qs��?��aNz�z��`���:*]�˘�xf��<[r�~^Sm�JKr��h����߼�Ƒ�t|`E>��$��Ag�)����j$��;&��7"�9�TBہ��#V��$�|.SK�ĠS́���F�_�����X�j�p#Ff�_N�(ϵi�Fc�b\�XР����ޛGvS��e/�S	D�D���V�4��7V�| ]j�i�|)
,OfK���)W"�xp���y-��5�
kպ���N���y.J�q\l�����n�%��Û{̈�ǃF�rnYvL���ЦC�dװ�d���G���h���<���3�.�L:�e�M  ��{�����y�хt����kJ�����/�$���i���aS3�Pٝ7�U�[zu��x�D�a=�`X>x�U�]L]��
�!�^�O��+��ǰ}�'��.����Ӿ�8���&�!4�,�ɼ�>xhӈ%��Y"�'Y�l)Dh��]�~�X�|��ۗf9�]{���Y�B��S��5������K�$�K����C��r��M?��$F��,,�$IS��NTx�o��`Q6�ܼ� ��cݚKD�S�%uJ��5����ʂ���-M�.�
�bx��=���$1x|3�����p�4�x���U-�ḧy�/Ҩ߉��oy�C��J}(� T#I�n�t����FRڷ�{�坏_(U�n�9DPZ+M5cb��\��dh��L�+ F)����.�6���_��nZ��*%q�,�K��f�&�R#B�3�IX���]��D@�ˇh�^�#��	$�L�%��	F�yD C�	��Tq�hWi��$�y�؟{�]�Z����~5��j����]F4]c2��\f���h̆W���w�UO��ԲB��љ(#�x
�m�Oa��0�G�sN8ŊU=�:T_Q�_oF�vżP&�0l���d՘&��6hQ
�-U�����4�a*+��U�FRU6m�{䶈�����oSAf��Ͼ@?��~��X��li:VHX굃uVmIA?c��1�%g�l�|^z 3�g�T��W
�,EM��F:��E�c;�2��2̡:+�v<Y�L���X�y�-��E��ь4N�o�Ft"?�M�ݑ�0��茨mWGc�L�f%��F���W�8�ׅ�oc����~��	��L��A��}���ѻO�C����4��Ի�����Di>���k�
��f���������X:QF���3ß��&�cTE'�ɰ�L�w����P�)���
�ף�|I�
�v$-q�kz��r�yLT���)	w�g�W�ƴ���h-X�H�X����;�����6��U�R2q@;����]�H�V�iNLP��K�'�F�<��Gn:���B����i2�_�'Hm����� ��X3{��o0"��:�ƙ�V�a�R��C{��^ߔ�����>o�\l�n��R2g'���t�0�?.���A��g=J��ul�m՛�i�W
W��$��V�&.�7_���� \�P��}�=;�O��N��|]?N���kH_��g0q.0��"멹o�sm<2�5H��Z����u���r�'%FOyv���ӕ�� �WSC�K_3�A��=]7V.�UQ �93{��bq���,�1z���y�b�b%�U��w�h0[��!���j^s�����1kOϊ�ƍYY�f��6�Z	2�t�#���D���;e4��2J���p�Af0	d��#Hm��M���}�5<�l������屚H��������e�:d}�E���MB���Γ�9����Os��A���#�Е�xot#�#nÇ�XS�҃^��
�ظ�`$*�S�'���,0��6����c���8���,�W'��Me�#M�&Lf�5��7&��DsY�����'H8�aC%��K���UI�w���Y0l�U}��ݗ�16&RQP����Y	LN�Ѱ:G?g��ʏ{��� ��n_zn��Er�?T�U��.�Hr4c�B�'pz{��3Ly��pS�����iK�O���8�״wRV͇G����<�݊fL�y�1=9��+T��n���ej��>������mI=ٷ�����$�+1 7�	�Ήǫ���t����ض�ob��t�;���|��ٷ���T�W=P����[$��H����/��"�/�MĴv�y��2�́}v�C)�6)qp$՗���帻�!��@A��
{}��!f�n�-�����)s�q�Y�����������.��weG���m�/@s�+�]B��� Y�u��&x5ic�S��?�U�;`MS�)�T�0P�z"�g7�c,�G�}��*-QY�z(��_�h���o�� &f�VR�+���ǹ��(�
5�A�̲�a����/����J�����ʗ��f�b�}P�BH��%�[v��J��E6�����b��$��訩<|�̱���w�`�]�
���Vƺ�W��7��y<.�KƎ�ǲJ/��$)��\r���VpDd8H�~���_��K�54��u���%\�L�A���}q�g1ං�'y�qd#�ݥ[^	�{�'��)�2�G�e��t�(n[K�	8K^�o
�*�EQ��s��-��a�K� ���;�gpӗO0��/~��X�[}{]b��(�k� ç�s��q�r��ʱp��is��R@�k�g5�Ŧ�Y(ط%�Re�G^�@��!%֛�zl��7���B܊�7M?ڣ�O��h�"�=���(�@ӟKG���
=��KEJL�*�a2�
�E|9��[��*ڝ����}�f%:���I|�֕Ȓ}t��g�^抱�^H�hl`YP߄��! g�RJ�LN�z`!!���y����~�� ��c���t����@Sp��UF��ʩ��U���*��-��By7�2��P'q7��+���rC����GMdx0��Y�n�r�C_j��ǡ�Ų����s����7�ހ"����̦Wl`�9R6�4��tO��l�_���N�K�X蜵(���Z@4�����e}v��,�����VB���.z���iw`���P�у� >M����'�O�P/��RĲ��M�R	kO�q�mYly76�xp��(:�ez��FX�{�1A%��OLB�E��$2��<#�$�]� ��6��֢(�ZR�/W"��e�r�������4���d��E���k�o�r+ⶓA���e���cu�(�>}Ҵe�j��� } i�����j�Y���V!�0�Qq��0���=�D��"�� �˅��p�ѡ��U�J�!P��:��9n�R\��anK(�	��*>�(�����}D練V��Rm
aY�-Bt'r�9X����}>Z�� �1�Ou��H	��i�i#7�]�u@��c��� �7�]�f�wE爝������#��zs:ä��)��m���Jp�;J:��|'Kd59y*���������B2����7*׷�fn�ݘ��	y�+Q/�O�ܔ�)ץ������ǒ���X33<Ԟ�M�����e>��n��$?�X��������So�z�m�61�X;}JlϤdiw�j������k9�2������cG� `������A�D���D����I�؆V&�3��w�m�v;��m:əy�x�wjc�O`��O�c����n'��0�B�7�^��%!!2Rx�f��f�� �8�U��R��x�}h��lO�]+��H��&�G��N �*�������@���ׯ�W�6b�����1ЗZ's�U!�>@5 m;����"ϼ�VX
�e�'g����?7���NC�x��_�&j4�J�O���WF��g&��(�\���x����l���� dRֆ��D*�*��Z��|�k��5I�ZO���jA'��E<� �Hwœ���N���j����NKQ�"�Gqei��Haq>3���>��K!&02pUg���bWE�3 jYG��]�nn�[),�QV}Vܜ�|�<��Wהv�?$`�u���dK���̛�Y�UhO2[S���Og
�&v��B�0r�F&S�>��䓤J(���cz���.���Aw����G(�� �_�s��s2�9�*�}���"�蜃�duhZp;J\`Y2���,7�h�C����^���=�+eNI�cq �^[��gA�I:�A��:�c6�RFбI��-����˅�����Z0�M��V�3��h�i�#��bu�hd���Å��!�F���Z�=��QE�����Y�{�(IC�]r�DY�/.<
&@����H��O�ꢀ�>�-��߱C ��co]x��{�:��??��/�p�E`�T�����Ks�s?S��R������G ��r�fXC�����q��M��N�h���]}�b��prvM�� �����_��Y4S��t�\ۃ�,1\(f0��L�*�P��Dہ�
����%A6,P9K�ة'5��-`(R���^.�nܦ+`��xrn�מ�GWA������/�Ŧ�ڲ�]��
{����g�}�{!w���Ӯ��D�_���=��q��?B����e�fJPb�D�P'%U�ל�R�cs�P)��|�:6��Щ�z�W��=��:N[2�ӡ	o�o&�2�7�Z-��1�b
�͋�$����	6�e�6�<�V&,^�0	��X'`$�tڇ�܉F�)�&!��z�6_2 .A]��I�� ��z���ܹ#�)����sV)��ν�Y^W����F�؅w�Y1��>���uݽU�!��UF�~r�Vߕg��B>��$�/8�RhaM�W��lFЎ���v;U��9�[e�z��JJ{�S��&�(I��,z��?�5�v�H�%��e�P�\d�[���WJ]t˝Y�염Տɮ�E>^� u�LT^�:�M��lT�K�V�F\j���-}W)(�~��:�/�;
�} �� ����kTU-�.y�(�׺��e��p�e����Q�ʙF[9p��Tri�_s�'}�tw��֬�8βCJ��َ�Fu���^>�qVAT�Ŵx�R�^�RjPZ 쯒�ÈP@'�`�}�8�y
p�I���B*������r8V�3QF��l����])�4~e�Cm;��9`k6Qw�Er���e�f)��:3@k��Y,����G�K�	�px��	a�P���Gb��B��f��|Ǭ��#1V�jڣ�G����64�a�v��C�7l��&A���>�F���B9-�ê~��`ně�����HK��/w2P����h��;�OCh�]UO�q��,��
 ���ȓ-|�p1#g!E�C����O	8t��U�{��r�e�m��s�+���@�oP�����'�@1=�(_�l1)���˦�!���teZ6�hTz]�F>�f��?�f��� �[�-���B��� }�\dq�)c*)�o+2����s��kaH p��3�e���\7xS�AȻp����8>�f:�? ������n37['gN�=�N;�/���P)��{�`ТZ=b\dù^�����_Ql�� ������!���F6g�p��e�õ��9mr����н�L#�!k�D�ֵN���X��8��H(@8�q�f����^��֤	zԌI�	ffg��s�<���Ec�p�YL�q/p�7fX�LAb�?e'p����ަ��dZ	=�+7qc�o���v���vG�����zT���I�\�n���l��`��td�S\�����Te�/3�-�Mdx�	)'BJ�4D6:$��.�NQxE�a6� S�0n~�)`������4w�D�r�2�|v���gE�R0&���c;���4��NV],�~�oR9g�"Ī��'ĩ����^�mb���)�GÃ�7Ϝ3מ�Sj6]�ݿW	
i��d���;�s�^�]�t�@yOC�	M��s�I����/�Ҷ���hB��mA<�L|��u�nj>�I��0l�ь�7�.�?d6H�y����s�x~��˟�1_[�UTB�e�_�#u�ƒ�,�D�8M�j�z����wG�@�̈�ŌpV�J�Ǟ��P�����euK����������e����'-�ί]Wh��ɲ�k2���H���A�T�VTR��x%.���;z-x��F��bW��]tǸD���6����Lrߚ����6@jG;|U���^���Ӳ?N�oX�,�I�&�h��.��������?5��Ǻ �|�\���x��+��Z�h����i\��#�Rg8�+w5+B��hr�̲ǿ������R�vv�bt�3��2/�M��h�`�Ep�mw�����Tn�O6|#�3�Q]��*U����}��kd/G����ȹ��]���F�w4Z/�12O5gZJ�\������oX�9�g�� ��Z{���O�U��%�*����7= ��J��{�����ɑ�y�����������R{�ݖ�I�%�a݈�FzA_li�(A��Y�8�@�\F2v��]�.G��P�u��Ⱅ��J5VN�t� AӐ�T4�|jA3��d"�Gѧ-��޿i2VKΒ�۔ȼ�U�D�1Tk�d�ŧ��P�Q3�R̴_�]9W���t�H�O0?q5g�NQe��k9D�6-�
j
�=�����\��Fnڦ�8z8���U!�؇q�5[��\m��0�B�,g�Lc��W-m+c�VX�������2�e-Rv���m4��D{"���k�v#�NLG�K^!�Q��J�7�������b�Jy�"�� ��g)��<+%r%ɿI�b$I��DMlNF��:h���|`��r��a���W)r���׌߽�*M�P�z���6�2�x��	�%Ѳ^�FLT)?��%�eq��ZAl�w}ؔv_�[ť���\D�}�g�\���1������=+Ɠ�V����$	�������A�%#���,6���+���Ռ�<��tn�L#��Q~E����l������p�dT����VS��}r��
��k�[���Ğ+����]����tyz�;�]�=���!�/߃<_NvJ��"�v6_�M�A��n�S� ��F����dj�y���*��;D��V4z��c��/K�.]�Wn��H��GW$;�V˕�2n��%a_e9 �f�ym.� ���y��7����z�ck��V8n�G?P7��<iV�EQ�I���c���զ 8+6�+��ѯ\)�uh�ܗ�ۓm��#�~!���Q���4s�Ґ���]�<���;X[�*t}
o���.��3�&��S{���Q��9��b����]%�w�j����	@!
VA�>RozLqHP���3�j�>���D�`�fHcS\��X]�{��+e�2T��A��E�t>�Pd# ��%d���45y�ч� z5<��ޟ��mK��O�?����$��%Ә
��y�4�'���F�]�Fw�?k ��
�/��s9Π`e�R���m}�=˷Em��"��ѩsW�.yJ��S�;��+������P�b��>�s��L|���kh�����W���4 ����fˮ�r��F�)Y� ľU��=j��j�^���z�f����V6u����.�i�j-T�;���ƇBiG�NM=!�������JM�]|1赟�ꞎ�[j�C�Ƽ�p�;{�Ϡ,l2a����TH�������ɚ .8��f�����;^S9�ʹ�S���ړB�Mg$��s���ʩ2�R�������:Tw㙈52������od�v%�#�#g;�Fw8�K�x`hE\�4n�&���8��I�&������
�U�O�FA�d��1O�| ��Sl8\%�����B�		�)�GUf5.B��Һ0�,�z[���I����p���VXIl�� bY���6 ����'�
{.׊��3`�2C:9�����}�EC�aߛd��h�Lk&%��"�[�P��fV��3��B��iڈB�u��Ш��g�mܔ��cU�z�]?��0��3�0��jۊk��<�ΰ[1�?���T�	��=��X\۴�:Q�(���PX�Qi�9�mN�/0��Ȯ�)�}���������_
m��^M\�Jه�R�4� �nl��x���F����t��qK�* A!T�M��D���$C}���
ypް��,FL-���:���0щ7�V�B�B	�I�kF��ub6��5����Ώ\��`T�_��M���V�sl�G��[�c֊��Ҫ+/�
ʓ8��n	#�O�`�~�s$!!�����X�RA8ߍX�,�
�B�jÒ]�*e���ǧY܋��rֆ"�Ʒ5~��@�|�j��3#�YYN�нe�'�T��Á�e^D�}��wwz[)C٦�2M꾶�����N�H_��/���Q���uF2ئUZ1;�AU���E���d����,W Ćc������K7 o��Q���>�W��o1\6�&�Ѕ��.����`���P�ͬ��f�Ж���x�\��y�l5�x�|@�'��L+|�,I�r&Ь�tg����p �U��|������v@�^������|�-�w��]�a)�5���E�P�fxUeeo��"�S`�ב~&��L'6�|����_5�wc�S	����1��o�ic����K�o}�$D��?�Rc�����/׽bS�f�i?�C3��KC�&����.���-�����[>�խ�a���>G�8�`�y�����Ov&��ۏ{����x��!�[y�s�k��Dj�/���k%[_x�dku��OB&��*P���sw��yj�0�@Af�+���E
e�X��$�.  ���-�'f�"�89�E2m8�x�ǰ?�
 ���R�O���@<h~�w�f���;a��X�i����(�Z�13���P��0��~"�dz�p�� �d�Ɣh�
�ɟl�p��I�D�9�U�5��'���\�Zk\���=Ӹ뉕����q�ٜ�Hu�ǀ�-ybY��
z_�ms�de�Ŝ!8���7��Bm��L��uU��?��ѽyP���������/d��@�Z1y���b�R����2(p�C@ꅧz���<@i�sf~���*��`�yE��,��Gp{���n�,ҷ��[��lͯ8��fF��&�O�]�R���߲����`i��O6"J6��GB�5�WZ����9c�Z-Rʹ���߲���Jobl$��3���|�<�����Q�*��<j�Z�GMqۄ�&C紙&XP���|D�
�:Y;�t*��`7[�ŀ�T49�"�-��#�x�d��0���'�|�?
&� �]T���������'�O9��+h�|�b���C�gG��c�-ME�w2�-d���7�R��y$*R��<]ﺝ!�S���k�P|ܬ��s^��>�e!�=|�-�f3�c�v��xi���9��$R��b����݅�
T./���
t��6�1bx�et��������Mr��.�d���/}�"�Yhr/����6�y��wv5@
��~��Ơ��;:{��R��lK���䭤0��'��an8VeL� ���G���twdv�-��Js�%�钲;O!�X�2*j���J��>�f[��G�>�B�Z�'�X��9���Y�Ӳ��]sZ�3,]����� � [�/lJpR�#������N+]�,~���ӓ*-���˥3�4��n�K-���bj�������^�h�����4�������E���m(��kP�Y�'����m����O�o]��QR�r�%���٭]on�Xvv��'������b-|@���d$��M
�s���b&ל�qEh!:��R�~�-��[�������l��z�G�<���K�e��G�F夆	?�-��cS_�w�QU��[y%�V�?�i�c0�˔r��}׽q�hK��J��YQ'U�O��f��.�ch�g���
NT��g'�KM��X��ж�p��l�4EᖭI��)�L`ٌ��GH~H(�_C��	���j}�J8|YT���S�aq�هN�Oq��o�F�����]R������jx���_4�C*��(�Y֌J�.�n	�,8Ӱ�?%p�ʏ��&��������@�<@��8��b7y�t��,�-�8>��VE�^�M�]����Z��i�<��"�g��w�����-��fqpʏNC^�'Z�E��efk���L�����Մ ˘���N�
*µ�#I�9��C]�D ��>��,)���5�(W{+}$tZ>�&|�g�����М� 0NrxC��Gd�2�n���ψ��1��g
G�\��J-Y���V{/+����h
�i&p��e.�d�O.�"gQ.�	B}H��U�P��Z#}�*D^�5��Yo�[�$�^-\ǿ���KZ�y����dyS0BwۀnXt�Nf�	��I�F��42�z8c7g7A���ͱ�	�E�_�U-�ˊ��u��8���.ab�3�ENa�=iR1�����4��[w�.��2���f�㏀A�OS1������eQ0�D��7f���h˾�"zg.#HwR �⨢�����T�#�΁�������z���V����̖|^�q��l�b�d~\�6�.К���>����e��x�z�)��e!pH:��X�aT��.���w)eʭ�
���K)W+�Q6�E�A�M�S�P(|�e�M�h�A���5�hW�C��@vY��MTJJ��"E`�X�F��Z���N���~X�P$[�Π;j�)�|�&�4�uP��~Ҳ�i��v6����7^<x�M& �d-�>�;���ɼ�+NM�1���H�y6�qT�cz��Ϙ`��i z��� )_*F�l:���'oa�
�f]����F>!o0���%���_ʍ&����$Z��|�}0i��"��+2M��KVw��=�%hr&�U�@T{�'��n��Ih*+��,�ʴp$Jۦ7HH�ݿ����K�Ev�K6����>��Ry8@����w�f�,���Į��U�V���5%�1���;N8�-�D����YP&}]�v��� *�m����K{|X����@)<��W�l�⾒�5퀮Z]���.���N5��q$��~R���4�cg�\���M��-o�-d�&��z���9��S�M����lyy�y�b����a;A �)w�J	bG��`�4J�]���
�Õd	h�����i��C�W�W�x^)+ X�+�_ �}�$z�`�y��:Q/^��af��р*���5'�b��$���W޺��C�+�
��
E���%u�ɳ�}��q��l<�B�W�Z;�b)�3ڟR�	�>��*��}����?�s�)Ʌ������NG\+dٜh�A���52g͝z?Q�gfvm���W��w�b�(`�{J�"*t�*���>�He���}m��$^�wH�ַ�Brg'jF:ǈ�	�?D�����?��a^�
�d�L��3��`�^c��+?ɶ�u6��į���z��+�e�}LC�N�ܥ�6��\hB���ӯ�&�<�#���E�;$���k��Ț�EG=����%:� �1�ݭ��ȐW�֯�|���YV��8� K0/��DHʀH�v!:�~I��09X���7��t�8��&\�#��鍯�0k��{�J(���sI�i��p</�'�����"���_�*�ha�K�gS�Q�d�����܁�0�(��OO�!Z%�������ϧ��,顉6m����Dxj��;��HZ87�
!�,3C�|TeNn�@*tgx&�#�	��dBZ<�<nL�.�n x�H̑�v�;��W��c�/�~�{X�]��ǝ	���7:[�5O-|�!kbH�t��ز�g�ӎ��#"���T�*��>W�W"\L��ـ@FJ�4����R��l�J�l��hi�1@�����3���}���K|�c�t�;�Ha�I�HA۲C�=����$m5ݔU�4�ٍ/&�ie�+�  ��W���j��uV�@���ŏ���=�4:�9Դ�OԺ )]ǳ��)_�1 �]��{l�3gݒJ��^�k��:��H�^1�n�����Φh�m���o^M��z)C��0��b�"������42��[�n)�ڧ��m���T\��X�3���C�x�7-O��uTa^��m�Ըޅ�:$�cczBK���F��\?ʃy���O��$!:����w��씲Q��i/���΄�}���64Et1��uI�	;��vlh�(C�3����r��v�����昀]I���������� o�KJd0|��ée���ӊ��=g6�Mu��IH�����\>�t���bFR2���V�`t��R��v��K�3N�*��Z�*��p�`wR��(G��n%"���Y_��Y#�S��0W1á�^����3Xt�y�q���B̏�B �墱k1:��e�2��l;������������c�EG�&���p37��}�@�0�v}
�%�x
,�ˑ����]�F̏�����$f�w�?�-�VX}O�1
�l	I1��(��N�9���I�A��ڌ���_�s<�� �n�!@�v��7Pa�/t�Dc�c3�����>���n6�y<�ǀ�6�E���!#�A0��[�E�?�ru��f[�р�ٻ,|���k�b���J0�~Ť;��"���&X���'?��f����ͽ��rf��ic����	��]��U��YC|Az(�	� +�� #���<w�ԿsY���R^4�y(����f��_]6y?���\�3{�,��!���E�EXD�{�[�?��0�P���D<��_��,��6� ��o0;�� g0>I��7J���?�Y�3���Z���rc�=�>au7����lZ�--W��\�$O�c7�Q����X��`�m����om_�^�Ы P;��~�J��� l�e�7�����u����I�ن7���H�a�*ޮ�r�ˏ��)����֜����v<�Ù��@�p'�M��Uέ#g��]3�����&<�W��J�_E$��7O_T&eg�ڬ3jU��EI��zсZ�,��żv��-��E@_�\a�����T�)h:E͗r駶�hlErh9��,���׿SB�?����_����y�7��r�v��[����^?�W*f����$.���T]G��p���z5J$�;��XBD��ⱋ�+b�-�Ǹi4�J�$9��]s�Z�5[�ב�A{(���	.#�c��Z���a�c������Jx[]}��!��#��������Z�C����2�m�RBX'B��s_�~�w���).'q����dQ����H�Nr��3R��/�.C���������j�*߶�������F/<9	u�":�N�/���m�iO�Ylw�6M���jQ��פ���U���jc�2U�I�9�x[��6�mƹc�1LFH�yK!�=�s�V~d��F^���{���_�a�1&��9�r���0(�ka
���1��9J�ܨ����`�I,/�%_x�ͯ���G�Z� Z�[LL�go�Q�p���\�y~C�,|~�",�1����tguD*�YfG��f%�@]�"ˤu}�� BM��6�K���6�!t%�'��b��w����r��~�~pr�������C��l4	�^>T�'E	Sg?�V�x��9I⽸������,%�!$���cx�X��A���}����=�f���D"�1W�����w�0�C�q�#�����ˠ��<�;�����F���qlN��L��2x?�� H���F��q��-��������k�7���{��QB�F�a�j�����7�D0t�%P��^�'����z��d�g��s���X� ��#�tFR7��I��u�7�9�39: ��`�	h!蟟G���d¯al"�l�?f��u�H?4���;7��8�� ��rGʹ�MW�(��R\�Jk�1��@Ĵ�m��Lu�#���nL	�ɾ#�O��	��X^h�>j�4/��!��.?_���>����PPJ�t݌^H��+w�@�m��f#H;���/x��HN��Bc�f�=R�X��.�����!<砤�Ń���i��ʒ3RP,�x��+��fk,X��|*��@��+�H��fF��y�G��u�3�7+]�hslsr#P�h�OU�лQ�����3�к���Z������OZo�r0i�������@L>����
�d�s�D���;�;RޔPL�����&8�l���'�jA8�#�+v��%:�3����?���o<LCxߢ�X%$W�Z��k�>"8����XP�R�f {�����k^�<� �&�B�V7�h\�
�y��e���|7X�$��d�=YU/�x�U�n�z!��NpM����`PP|�r����69���q��}�Y\�Ɩ{��4@���j�n����n�ճ:�A3���#$4����;|�-��s�= G�Vx-���%"e���Xo/��d�����?v�k��Z���LL,��qKp�����ĐQ�Kq��qt�� ����.c9)1�\�޹�R�:p��)�g�߮ѽ����n�����R,�IN�:#�TY��^
q�0�� ��yD�	_4�[k:Q�R�`�}~v�ץr�u�ܟX����r��CkV)�y��Ҹ�t�I���|�^J��X�}���������V���%�q�`�:FI�Mo��xv�,��܈$<Kc����+W8	�fJ��uZ�UvZ�*:�Ft�'48J4C���V��Knz�����3��y�h���.l�r����%S��G-�i���H�f��p*����n��ᡨ_>��u���]
OrP������Z�`�h�!��q�j�#��������	<e��ҿ�!���5m�]�
=Y�����G�Ȗ�<�[,���e�;nH��ǀ��	�7��T��0�|���YR��Vx7�v��I����PO�x����N���ki%�z_J��x3�+��Cq:�-�xKP	�N˗��8ΐ �}*�m��ܠ6R�P�_�)�1s])����tdF���;�"�$�1bt�]Qw�tT���quL��ih�O��r��/\&F)�D����ʾR���87��<�� ��]f|}E�+R/�I&�^�>�"ȍ�I͒���s���a����| �� o�"��&�R���?*?�O�A>v�jlq(H@|.c3X�HL� y�m����hǧ\�����ׂj]Er)�+Ii~I��+���#i]|�:kD+@�7q�.{��Z���ׯ����Gm:�<� �K�����V��8�Ŗ�Q���V���6���x`K,�ot�s�_����2�=�fW#҇�:��W���Y	��+˾��$���\�S��e�p�i(a��+� �Z�>���U=tPn������_<iOۮl���X!؅ɪ�q=U��%���t�c3��&?&<��Zy��� 7-+��Ս��G�(]�|�����R�|x�����O$~eV�G���{\�	<�_M#jk8c��QQ����BL�D����-��*ͮ�J''��
�b�v*Hi�-<i��no����f*�Yb��W����mۛx5}����m���'A�|9Y)Ww)�0Z�40�:��N����Q�u��^����L�Hl��ú�rn�����n�o�n ��3�;�'�H!�;�^��Lܽ��%�0�M�v�"�.�) ���x<�RTaɏ��#��᫔��st�*y��ۏ�[�|&y�+{�{c���C\z"	��v2���6:�BN�E0-�&z��ݧ�D��Yp�g#�6)^�q�6@�)s"H��r�����&��G/��W�Uʙao"Tǭ��LD˂�W���'��=��[���r
~&��a�Iu)�	����-���'!��͟�[�`���Y�s�9<�dxX�^����v���*�1S��l���w��c?N4R}wg�̓����E��`��t��N�N��"F���#,�L{��	����5G������3�����3F`$����9�J�en�b���0�W��-��֬�gv�.SҞ-�D�*2���qe������o�~jo�m'��eò[)��|��K�����5���_`�53�lWu�vj�|���T��H��7��r��o-t��ʀ�q�Y�<�N�Z����|ŎK߲��ע��ӅK�c��=�\׿���7��`�U[�tqfuZ�����.
*��?9}/��<@��6�79o�St���-� ��xo��^\}G8T˩�����}�g����-N	�Le�1%�W��Qp�$���*���-�똱A�w�G��(�06�3�r��-����LA���м�O�z]Ld�F�3w�ӽH$g�L� ���F<�$�~,�KQ���~��ŉ�eH���)A�hs-�6IU60{�ua�:.�hшtw����$�!b�u�9�V����n�(���(��w���i��]x��[��S'e�g��������ȇ�an�iAB��������چ������^���!�ю��]F]i�8��?z��B{�uY!J��KQ�T���av��5��+]r&��J�[���\�r��j�y���K�f��p���>г��o<�_(x��s��� ���k��Ḫ��{"�^���?�����/g����V9&f�(�mv/�A�n���\�S��r� !(+p(�C]���֌�u� �����-r�x��^�6������qc��#N'E�aCxޔ��E�h
�N?Z�`����2���QԘ�(�w_��?دVcz�.�\ܣ��F�L��9
؛��]�G�ɂ��`H�^���o��eV�V-�}��|��x�p�l�����h��˛mc����,q0qy�b�*��yԗq�UI9NC�(��<-�@cZ����xJ^Yz��USr$%�
&���~�mEe�L����&�)�7��<V�+{QZƻ�0_���_eg��������:�)��a�Y���$z\���'��_f��n{�8�R��1��)_%'˒�ץ��G1#��Z����v�����8��	��Pn1m����Jz�������H"��~�vICS�5V+��X��9l�dJ��է�������?S��Ub���:Ίa�b����^�./�&P'���P.s.z�q���Oq�d$�z���[y�"����N���T�h+�-e�H���DC\��΃���%�vt3�[_�N�d���)����C���,6)����U���x}p���xw��uTT���p'[�m+U��y�+�-���o�<�j���7d�
���-�>m	�Z���r�p��kc���YKmG���y~Njڧp����y�s� ,����t�dS�b���wt:J=�ƚ��ʍ�g��}�H�бԢM)�͞7F?��h���[ɵy���^����vȧ���)5����`mh0��a2��_���3*��U6/�z�(n��XR</��-F�K��܃��ѐF�8J������jS��m�C��2��5z��4�deM{�·6#d:;K4Q-�\�\S��O����ܵ4ƌ�%�
��ٿ~0�u���˄p=��巓�l��n�?�,xf�蟄@�+��$Xu(����U��'c:����\^#��;3�0�\D/�0�"�P�,�V��������Nr~LUbڻ��=-x���]!K��t(V�6�N-&�����бF8;�	oD_R3����*J��R�rWya5j"Y1n
Y�/y�As�l۱n��v��ݵ�~�P�\o��u�PJt��ɉJ���X�.���Ei��$Ym;�����TRi��g`��L��+�#gH�Δ����?G�j�������8��/��=މ�����@Ղy`H���<)޽ݟhl)d�kz2����wP�Fw�.1�&�|�s�eZ��,%l�J4���w��@���g�i�-K�_�D2k��I9PMn�ʄBI/��jYd[/�Fi ���)��*"1K/�p`�ߥ�*�C� r��M����E�+�����@k�H��s���+�Dg�ߑ^��*]~�ܕXV��B;�[ǁx�B�ź`��3,�`,�p%o�.o���jvd��r�� ��o1r�0I@wF�)���:�R+� ����c�'0=C����edU~,���Ϗ�.�eF�Ӊ0��Ӧw���o��v�����a1���G)�̒��� Lb����(�(V�zE��i	�����66�!�:ܕ���G�1����Zֿ�eدyy����ʈ�$Q�'$l�x��,�ka��H�����^H�4�L���WdS��k��
��9ņêi�ӿƭ�����m���D��wSzh�p^���;����9�?l(��Y��8y{�����������T�����A0M{�[�ܧ���
���g�FRͫi�7	��	=��ߊ�w
��9�*8\*~�6�ܶД!(X9Qǭzv����~�85q�E�3Ʀ�G�S�1�M�S�� Z���MX�~���nӏ���~�NTfZvnp8��YEx���h�8TCVJ�#���k*�����B�,>�M�Z�ףF���m>r�]��P�K��t�m�`'����#�%��~jWo_+4U<�%��0"D�1s�6�<5��t��:+�w����sH0�A=Y�ܹ$V��)�f-8R-�28���J��*x�l�b��g����#!>��K���鱴��w�{��A�bzQ�k�;|ϚgM(ݙ���JƦ��726�Ww�hA��51q�K3>�R�"�I&���D�I##g�в�cq��d9��E &�tgǐۖ��G�����;E�[���a_%2>�.��:u���2��`tv�F b�sA���I�_سx؅�)gK��,b~��t��X�R��{��?��J�#_j��C�i����G8��J#4�F�+t^�r\���v��$�$����ןc�!������#�N�p�b�~|���=�u�m����k��Ÿ�pN>U?wx^
�$�{L��Y����W����?~_�qMl���ȭX��t�������e,��y2)�K9���gC�����	��@������Z��8��c��5��
AQS��:�A�d�ʯݎ,�{2Hn�ks�I)�κ�ɵ�0��l��h�7Kc��<j�5ؖ&��+�-�pE˕����m%���u��r��ψ�B���5�d��]?�3-�W�f��0s=RR��i怜+��w�D�M�X�r�����%&�ؤ���KΪX�֛6�.!{��&=�>���ěH�@Ū�U!z��Q	0|�$����!��Q��}(6�L�Onİ9Um�;�A�4x�T!�F�EB�~;������J���*IL�1��]��?2��W��!r�8S�@�1L;$�ɚ�2S����kTE�k�@�(�Z	[Ŷcya��e�9:�yŸ��'q$����6�e��n0Y�!����So����>4F����B=���Ua_��l��o�^�cj��a
�#�sQ@y���;�[3y$>���A��tJ��qܻ;��Dc
�8�B���͛���	Մ��K��ϏH���ω��Y���1�-��t�y�[%M'�a����3�����mx�;�k]����n>���yDA.���Scy�U��1X�|E�����:b�^� �юaZ����S��(���^�*�~�K��F-Z���v�3Z,�`���?���n>�_&�?_U�=g�2�|�s��R�KX�-r睶#-����fZhi��Y��_s��Y3џ�+��l��B���~��E20�\E�X�[���r.��IX��$��?Y�Ө��ɡ��25��o��g� �����ѯ�kڶ��R��8��0mܜ �=|��%F�g^l�ͫ1}��n:i��E��cl��첍Z��itPJ'�d����������a���&�7��8�1�ro����"��I(@��g�"��]�vW5?Vm#��D�\����	�#��2O)\=���.Go���Obl�y���%��n����N�XE��e�D	�>Y��:啝?�F�>an��}�ߞM�v ��5��7�e��`����Y�b�4���ࡒ<�B9 ��R ��$� G0�Q���� R�)���O�%M9��I��ʄ�7v�$�D� RIA{�k{_����C�OM�/�u��>_)��m���N�![��7������hz���&Rfxa~ɽ��]�h�v,h��vD�Es���9��%P�mӟ����l��95��M��ؗ��$:M.����
j�9����ͫ^'�$�ݸ��7���j�˻���׍l��0I��C<X��,输�	���_�Q&*D.C���{}����H�baވ�Ϛ%�ak(\���Y��诙�2�^�=i~O�x��4�E'�O!����8�+Y}L,y���9����8���wKiZ��N�Z؁�j�BX��{���(��x��U;[7l�X��.�jQ(A�b�pD�{?�.6�:�_� �qz��i[\�+�v4�����9X�4��z��9���w]�y�n��A{UY��S�k=�����_R=m�	Zi�)����B%'�i�އa�,_*O��ә����)�[��_�%.y�".^}H ;m�f��xh�T_���!T�_\ #�αF[	3Q�Kˁ��~؉�$l��0ۓ!/B;��k��o�6�� Yg]	�/��j�%�r�~EX7:Y<x�m0�̕O�Kq3٬�K2��h���ğJi�z��(y���?��d�� � ��a����hJ�}o�Q� ��߯>cn�YB��X@r��c���1`{aa"��P%��Xlb=&��r�
%�v/�^����T��A#}����ry�E�c����ωL2u��hr�����#ዲ��!��C��M��T��茩�Ev�m+��n�W�������%�M�J'7Jv
�0�zE=E[�Fȡ���D/pI}& a��M���:��9?f����wm�E����l�>�Ӑ:<�ƿ�`#
�����ӛ.�=k�^شDF��M�GW�Y��\�\<�0W1Ή��G��nCQG؀�i��tP]��6S���dR:��G�'Ek�� oe�p(���G�c�z�����258�A����`�{i]^^�H�(����`�����]���4E���u�I�Ȱg��z[bA���dɚ����o04�#��3�C�;�@L�D����>o�\��ϼ,�,� �E��������䕿#�&+��0�jHWoi��}��0bH�i����`��R�0�@*K�dVQ�Ax�����gIP�ޕIQ�H
�x�iA�R�g)pt	�#j����N�.��x1c�1=[$3n2&Y����Z�%
��D�<yNLx��9	����_���rfK��Ҕ��ChJ��.3l��p� ]�|0UN&㫗{۫��q�k^Uu�M]�:�=h7ʍ��u ��ڸ��D�|e��n<F ��PS��jَ��K�a<���-j�>�r�| &!٘�,� >�7W�a�uC�f/�!p׀����/�\�K�9�ʑf�ĭ�c�}�c��Q��0{Ӧ7��G�+�#&ܕ%����Ag�H�.�I&t'��1�T2#x�}�Z�F'S'a�[�7�Yă�S��'�6�'$@��G�o���<l���sY���h̪iK���w�>/��IP��g���Βk���L�b��N�^����m�i�K{�X98G튧,�?�(�6���krW��Xj�}��� �F$5��B��I�7=��K�$�h�����%h\��q6���x��q�E�Ǭ�'X����.t+O���+ckXF8қ �B�{?����;�b+%>ۗ�s��;���~�����p͒}�ƾ]E�/8օ@j�	t��W��# ��U]��Ո�I�� ���LN̵�W
F��v�	��^������)P��q_d�(Z��J_�1*��n QBK:�J-�"���0�iũ.���B�Z�-ۖ�eJ���������7/}�����m��-��N͞	����g�⊅Sr���9"$㰻���Vm�c�B
�#�9�Ķ�S��/��ն�я%��1Mmέ,�<����͓[Nk�;Cي]9Lo�lT(��?{:�C��%+@��?��c�]��Y]�t�ɋ�,k��Q��o�C[,k*ܻ����6�Q޸��SaE;��m.f�"�Z�r\�Hm���$��K��q`˕z
�҈��.��_>h߬���<��l�QU���9������p�%r?3��9y E��j�0}6^�R_��LG����n�aFF��[����X6���VA��Fw��G�CX[;D��j3�����r�����5g�i��h�:F����tG���#Yx0����ke�{�l�W-@�9�@Lʥ�9ϕ������f���SaA~�@_�@�y���WԂ�Gc�9	.��P�F,^?N�V�������[�Х��ci��"0A��<�T��>�mvI}㓨�U��s�_�>Dj�`��s�~��c�v3����|&�I�v�4����>�f2��Aj�_�q��'��CD�~UG����
0O;m�`�_^��yd�B*��t��<��@Y,�ʋ��U�H��c�$���m���(J��_M}}Q9�6���Ldd���e�5��o�K2���{K�J���(G|��jtl���=���X���l�o����G8�`ηV�]�ڑo3/.�O�;I�v����}�+���&�^��ʺ�ӷ�ں��JzB}��&��S0�:��JU��媄�)�N¨�C�G����>�G0���(*x��PM��G�^v�ȿzԌ�3�6��%�#�Ъe�W�7�
�k3��gژ�7H\�J�����vI ���|3X3Ǯ��4�z޳�,:��V�������~��c�,�T���������\躒���}	����w�r��ۮ ���ۏ��T]D�Pw�:@<d7Q6VO�O,��0~ �e�:��m��|�O[�QRَl~��f�~��!/�������n���J����@�:��ûP\��=v�W��.Yai��1e���cO�O&fKY��)t�J�D}��>3/�2w7i���#QF����O�q"��;�Ӷ�8�/̙�����8�N��k�8�G�����PR��(�d-\��"n��}fT�3'�	G��6�0Rc�T�L��#����\�`T�`Ȧ�-!ӵ�<N#�@�436��-�.�2:�e��`R�a�5��,)>�?t�����-�|���� Y<x�m��r�������P3��o����+�O�v����l�<#�i�����;�vo���W�.�5h!T�Q�4�]k�R�	�K&So@W,����_ m��7r��:��4�d�ǧ��5�wo�q��{4�Z�H@Y�%,��KKE~d���aK�A$��t7nz�#�e�X���ew��� G��`������f�P���������~Z<�YX
�Y�F
�@0��c�y�W,nع�l}ʔ_gW��k��	��ֆ�0�)�[��W�yu>�����|�Ƿ���d�؜&G���P��;Y�Y�Pr<�gL~]�	�q�LղO�4�_�]��3�T�a��&~�ތ�R��9��e]�!gP4^V�����|�[���c�@�G��H���A����k$��я{�j�f
��� ��'�#6#�C����	8�6k��w��A#�˜��9y���+iasc*�v�l�H�A�M��Lq�����z$_@d�`�|K@u0��K^قypr��6����@�ݽ�<ڢv�3� ��O`��$�-�����pH��t�`b}^�̘07p���®]'�"M��R��.:�<���0y���lj�B���y�pPu#��S�����.�e�zR����,��Rh�f
/��}�}���&f#hE���%��T�)���h�P���-Ce���i�e�6�Uo�rT�;*z�K��X�x���!�C�/�Hl�%��pS�9��a,�H�ڡkdP�Dm.�!�{n�ҏ�<k��&�����B��!:F~���f��(`^������:��v-�}<`]Dݑ��,+�*;H���o�tl���WO�������| `����!�"��&��Ԇ��MO�DL��&QEA�Ȋ�j�B����Hz�" ��od�ԁ��E,eņ�Ĩe\oמR�g ���� ^Ӏ�4��ȀT苣�L��<��dԽ�U�c��SEl��	��ϰ>�y�W{�$W��Y�d9���Mj�9DsP�^����ME�J4K�[)ܯ��+75Sᱱ�u����8�hL�mC����1��������:��i_��2n�s@�� >��tNV�3{���(��}����Ӑ"��T�Ӎ^RV\>JfSӤ�cQ�z|��+9	y�c	?1�뙯e�,۵����L�uM	y��'nޠ�[8D��	���;=��[fҥ�yW�H͚r��-AV`�7a��vC�4pE{� ���\�D�L���'+�ٿצ�啴�;��	�q:̛�t;�Ma�$�7�K����a]w׵��9�a˔y��@��9���jGYy%�&aMmoDt� ��|)|KݍO"��bt\WK�G���W
��ػw���O(�!`��c�л���ě(�.��/n��]\:�s��)�P�Ի�_Cs��Ek�9ah%�"�OR����Q�,.�R&����sU�����2��!�UShsX�_:�1�N�v��LtB�p�^f�H]Y��s����QڰSUNY!C�#�Y�bf�><�;��i�I��.��MP�_�;����&5��!���� ����.�tȌ��<��$H�x�0s�q�v�t�IF�N p�a�s�0�#���ҮB+EC:�� ��U������=_M��:Ny�lG��~�Y�w��\�X*�+����qJsU���RTSA��SM=�٪�"o�рF�8�d�z6�d0��� 	�8����o �#�"�,�ra�&X�[[VXm��Oa�(]����λ�s7m�q�����ͬ�+]1��G��b���m̒�%�fOX�QLR����;�#q�c�<X$eW��g��u�5-���X�kbҥ���,lN;��4�H�ԫ��b/�L���YG��tH�'��ӓ_�'� �#
�:�)���\E�۸FD4�lvd�̝�����1k�����\��p�FƢ�Tj!ڰ��f��h���Q��veU%K�Җ�c�zs�Y5}k;d�q*���?,���?����"��׆���Uw��p�������(0�
�,�(SS�B�0]���l"W�~��e���(�2�Z��~�!�q�iG�ϖ56���=��F�V��ɬL�1t��+��b��R���� ��QUF�ǭq8� 31����ޣ�����c��������e;z@K\�%룸��k�8���q��koWP;���[�g�:k�EKB��h�k�o[���O2�I��珊�0�8�,q�C�pY;���{޹nBVIR��Rv�I�by��<c���*��3i�җ����������Tbo2V�8b|�_a�<�;Uh��s^%��
, ��si���`ë�R��r����8*Փ"�reȂ⇖9hg�	S_����-R�	A����E|��I�����2^fBD���4�(]VO��ݸ�9
/�Z,I�T��]�!-�A�XOh%�boJ0QXS�I����]��?J�}i��ڄz�+|�9���9l�X�(i��Q��\&��ɹ�@{���I