LIBRARY IEEE;

USE IEEE.std_logic_1164.ALL;

PACKAGE cos_data_pak IS

	-- Define data types array
	TYPE data_t_rec IS
		RECORD
      		data, result : std_logic_vector(31 DOWNTO 0);
		END RECORD;
	TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;
	
	-- Define actual data
	CONSTANT data : data_t := (
		(X"00000000", X"40000000"),
		(X"0066F196", X"3FFFAD35"),
		(X"00CDE32D", X"3FFEB4D5"),
		(X"0134D4C4", X"3FFD16E4"),
		(X"019BC65B", X"3FFAD364"),
		(X"0202B7F2", X"3FF7EA5D"),
		(X"0269A989", X"3FF45BD5"),
		(X"02D09B1F", X"3FF027D5"),
		(X"03378CB6", X"3FEB4E69"),
		(X"039E7E4D", X"3FE5CF9D"),
		(X"04056FE4", X"3FDFAB7F"),
		(X"046C617B", X"3FD8E220"),
		(X"04D35312", X"3FD17390"),
		(X"053A44A9", X"3FC95FE3"),
		(X"05A1363F", X"3FC0A72E"),
		(X"060827D6", X"3FB74987"),
		(X"066F196D", X"3FAD4707"),
		(X"06D60B04", X"3FA29FC8"),
		(X"073CFC9B", X"3F9753E4"),
		(X"07A3EE32", X"3F8B637A"),
		(X"080ADFC9", X"3F7ECEA9"),
		(X"0871D15F", X"3F71958F"),
		(X"08D8C2F6", X"3F63B851"),
		(X"093FB48D", X"3F553712"),
		(X"09A6A624", X"3F4611F7"),
		(X"0A0D97BB", X"3F364928"),
		(X"0A748952", X"3F25DCCD"),
		(X"0ADB7AE9", X"3F14CD11"),
		(X"0B426C7F", X"3F031A20"),
		(X"0BA95E16", X"3EF0C428"),
		(X"0C104FAD", X"3EDDCB58"),
		(X"0C774144", X"3ECA2FE1"),
		(X"0CDE32DB", X"3EB5F1F7"),
		(X"0D452472", X"3EA111CD"),
		(X"0DAC1608", X"3E8B8F99"),
		(X"0E13079F", X"3E756B94"),
		(X"0E79F936", X"3E5EA5F5"),
		(X"0EE0EACD", X"3E473EFA"),
		(X"0F47DC64", X"3E2F36DD"),
		(X"0FAECDFB", X"3E168DDD"),
		(X"1015BF92", X"3DFD443A"),
		(X"107CB128", X"3DE35A35"),
		(X"10E3A2BF", X"3DC8D011"),
		(X"114A9456", X"3DADA614"),
		(X"11B185ED", X"3D91DC82"),
		(X"12187784", X"3D7573A5"),
		(X"127F691B", X"3D586BC6"),
		(X"12E65AB2", X"3D3AC52F"),
		(X"134D4C48", X"3D1C802D"),
		(X"13B43DDF", X"3CFD9D10"),
		(X"141B2F76", X"3CDE1C26"),
		(X"1482210D", X"3CBDFDC1"),
		(X"14E912A4", X"3C9D4235"),
		(X"1550043B", X"3C7BE9D6"),
		(X"15B6F5D2", X"3C59F4FA"),
		(X"161DE768", X"3C3763F9"),
		(X"1684D8FF", X"3C14372C"),
		(X"16EBCA96", X"3BF06EEF"),
		(X"1752BC2D", X"3BCC0B9E"),
		(X"17B9ADC4", X"3BA70D98"),
		(X"18209F5B", X"3B81753B"),
		(X"188790F1", X"3B5B42EA"),
		(X"18EE8288", X"3B347707"),
		(X"1955741F", X"3B0D11F6"),
		(X"19BC65B6", X"3AE5141E"),
		(X"1A23574D", X"3ABC7DE5"),
		(X"1A8A48E4", X"3A934FB6"),
		(X"1AF13A7B", X"3A6989F9"),
		(X"1B582C11", X"3A3F2D1C"),
		(X"1BBF1DA8", X"3A14398D"),
		(X"1C260F3F", X"39E8AFB9"),
		(X"1C8D00D6", X"39BC9013"),
		(X"1CF3F26D", X"398FDB0B"),
		(X"1D5AE404", X"39629116"),
		(X"1DC1D59B", X"3934B2A9"),
		(X"1E28C731", X"3906403A"),
		(X"1E8FB8C8", X"38D73A42"),
		(X"1EF6AA5F", X"38A7A13A"),
		(X"1F5D9BF6", X"3877759E"),
		(X"1FC48D8D", X"3846B7EA"),
		(X"202B7F24", X"3815689D"),
		(X"209270BB", X"37E38835"),
		(X"20F96251", X"37B11733"),
		(X"216053E8", X"377E161C"),
		(X"21C7457F", X"374A8571"),
		(X"222E3716", X"371665BA"),
		(X"229528AD", X"36E1B77B"),
		(X"22FC1A44", X"36AC7B3F"),
		(X"23630BDA", X"3676B18F"),
		(X"23C9FD71", X"36405AF5"),
		(X"2430EF08", X"360977FE"),
		(X"2497E09F", X"35D20939"),
		(X"24FED236", X"359A0F35"),
		(X"2565C3CD", X"35618A82"),
		(X"25CCB564", X"35287BB3"),
		(X"2633A6FA", X"34EEE35C"),
		(X"269A9891", X"34B4C211"),
		(X"27018A28", X"347A1869"),
		(X"27687BBF", X"343EE6FC"),
		(X"27CF6D56", X"34032E62"),
		(X"28365EED", X"33C6EF37"),
		(X"289D5084", X"338A2A16"),
		(X"2904421A", X"334CDF9C"),
		(X"296B33B1", X"330F1068"),
		(X"29D22548", X"32D0BD1A"),
		(X"2A3916DF", X"3291E654"),
		(X"2AA00876", X"32528CB7"),
		(X"2B06FA0D", X"3212B0E8"),
		(X"2B6DEBA4", X"31D2538B"),
		(X"2BD4DD3A", X"31917548"),
		(X"2C3BCED1", X"315016C6"),
		(X"2CA2C068", X"310E38AF"),
		(X"2D09B1FF", X"30CBDBAC"),
		(X"2D70A396", X"3089006A"),
		(X"2DD7952D", X"3045A795"),
		(X"2E3E86C4", X"3001D1DC"),
		(X"2EA5785A", X"2FBD7FEE"),
		(X"2F0C69F1", X"2F78B27B"),
		(X"2F735B88", X"2F336A37"),
		(X"2FDA4D1F", X"2EEDA7D4"),
		(X"30413EB6", X"2EA76C07"),
		(X"30A8304D", X"2E60B785"),
		(X"310F21E3", X"2E198B06"),
		(X"3176137A", X"2DD1E741"),
		(X"31DD0511", X"2D89CCEF"),
		(X"3243F6A8", X"2D413CCC"),
		(X"32AAE83F", X"2CF83794"),
		(X"3311D9D6", X"2CAEBE02"),
		(X"3378CB6D", X"2C64D0D5"),
		(X"33DFBD03", X"2C1A70CD"),
		(X"3446AE9A", X"2BCF9EAA"),
		(X"34ADA031", X"2B845B2D"),
		(X"351491C8", X"2B38A719"),
		(X"357B835F", X"2AEC8332"),
		(X"35E274F6", X"2A9FF03D"),
		(X"3649668D", X"2A52EF00"),
		(X"36B05823", X"2A058042"),
		(X"371749BA", X"29B7A4CD"),
		(X"377E3B51", X"29695D68"),
		(X"37E52CE8", X"291AAADF"),
		(X"384C1E7F", X"28CB8DFD"),
		(X"38B31016", X"287C078F"),
		(X"391A01AD", X"282C1863"),
		(X"3980F343", X"27DBC147"),
		(X"39E7E4DA", X"278B030B"),
		(X"3A4ED671", X"2739DE81"),
		(X"3AB5C808", X"26E8547A"),
		(X"3B1CB99F", X"269665C9"),
		(X"3B83AB36", X"26441343"),
		(X"3BEA9CCC", X"25F15DBB"),
		(X"3C518E63", X"259E4608"),
		(X"3CB87FFA", X"254ACD02"),
		(X"3D1F7191", X"24F6F380"),
		(X"3D866328", X"24A2BA5A"),
		(X"3DED54BF", X"244E226C"),
		(X"3E544656", X"23F92C8F"),
		(X"3EBB37EC", X"23A3D9A0"),
		(X"3F222983", X"234E2A7B"),
		(X"3F891B1A", X"22F81FFE"),
		(X"3FF00CB1", X"22A1BB08"),
		(X"4056FE48", X"224AFC78"),
		(X"40BDEFDF", X"21F3E52E"),
		(X"4124E176", X"219C760D"),
		(X"418BD30C", X"2144AFF5"),
		(X"41F2C4A3", X"20EC93CB"),
		(X"4259B63A", X"20942272"),
		(X"42C0A7D1", X"203B5CCF"),
		(X"43279968", X"1FE243C7"),
		(X"438E8AFF", X"1F88D842"),
		(X"43F57C96", X"1F2F1B26"),
		(X"445C6E2C", X"1ED50D5C"),
		(X"44C35FC3", X"1E7AAFCD"),
		(X"452A515A", X"1E200362"),
		(X"459142F1", X"1DC50907"),
		(X"45F83488", X"1D69C1A5"),
		(X"465F261F", X"1D0E2E2B"),
		(X"46C617B5", X"1CB24F84"),
		(X"472D094C", X"1C56269E"),
		(X"4793FAE3", X"1BF9B468"),
		(X"47FAEC7A", X"1B9CF9D1"),
		(X"4861DE11", X"1B3FF7C9"),
		(X"48C8CFA8", X"1AE2AF40"),
		(X"492FC13F", X"1A852128"),
		(X"4996B2D5", X"1A274E72"),
		(X"49FDA46C", X"19C93813"),
		(X"4A649603", X"196ADEFC"),
		(X"4ACB879A", X"190C4422"),
		(X"4B327931", X"18AD687B"),
		(X"4B996AC8", X"184E4CFA"),
		(X"4C005C5F", X"17EEF297"),
		(X"4C674DF5", X"178F5A48"),
		(X"4CCE3F8C", X"172F8505"),
		(X"4D353123", X"16CF73C4"),
		(X"4D9C22BA", X"166F2780"),
		(X"4E031451", X"160EA130"),
		(X"4E6A05E8", X"15ADE1D0"),
		(X"4ED0F77F", X"154CEA58"),
		(X"4F37E915", X"14EBBBC5"),
		(X"4F9EDAAC", X"148A5710"),
		(X"5005CC43", X"1428BD38"),
		(X"506CBDDA", X"13C6EF37"),
		(X"50D3AF71", X"1364EE0B"),
		(X"513AA108", X"1302BAB1"),
		(X"51A1929F", X"12A05628"),
		(X"52088435", X"123DC16E"),
		(X"526F75CC", X"11DAFD83"),
		(X"52D66763", X"11780B65"),
		(X"533D58FA", X"1114EC14"),
		(X"53A44A91", X"10B1A092"),
		(X"540B3C28", X"104E29DF"),
		(X"54722DBE", X"0FEA88FD"),
		(X"54D91F55", X"0F86BEEC"),
		(X"554010EC", X"0F22CCB0"),
		(X"55A70283", X"0EBEB34B"),
		(X"560DF41A", X"0E5A73BF"),
		(X"5674E5B1", X"0DF60F11"),
		(X"56DBD748", X"0D918644"),
		(X"5742C8DE", X"0D2CDA5D"),
		(X"57A9BA75", X"0CC80C5E"),
		(X"5810AC0C", X"0C631D4E"),
		(X"58779DA3", X"0BFE0E32"),
		(X"58DE8F3A", X"0B98E00F"),
		(X"594580D1", X"0B3393EA"),
		(X"59AC7268", X"0ACE2ACA"),
		(X"5A1363FE", X"0A68A5B6"),
		(X"5A7A5595", X"0A0305B3"),
		(X"5AE1472C", X"099D4BCA"),
		(X"5B4838C3", X"09377900"),
		(X"5BAF2A5A", X"08D18E5E"),
		(X"5C161BF1", X"086B8CEA"),
		(X"5C7D0D88", X"080575AE"),
		(X"5CE3FF1E", X"079F49B1"),
		(X"5D4AF0B5", X"073909FC"),
		(X"5DB1E24C", X"06D2B797"),
		(X"5E18D3E3", X"066C538A"),
		(X"5E7FC57A", X"0605DEDF"),
		(X"5EE6B711", X"059F5AA0"),
		(X"5F4DA8A7", X"0538C7D4"),
		(X"5FB49A3E", X"04D22785"),
		(X"601B8BD5", X"046B7ABD"),
		(X"60827D6C", X"0404C286"),
		(X"60E96F03", X"039DFFEA"),
		(X"6150609A", X"033733F1"),
		(X"61B75231", X"02D05FA7"),
		(X"621E43C7", X"02698415"),
		(X"6285355E", X"0202A245"),
		(X"62EC26F5", X"019BBB42"),
		(X"6353188C", X"0134D016"),
		(X"63BA0A23", X"00CDE1CA"),
		(X"6420FBBA", X"0066F16A")
	);
END PACKAGE cos_data_pak;
