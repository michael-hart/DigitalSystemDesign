-- first_nios2_system.vhd

-- Generated using ACDS version 13.1 162 at 2016.03.04.17:29:02

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity first_nios2_system is
	port (
		clk_clk                            : in    std_logic                     := '0';             --                         clk.clk
		reset_reset_n                      : in    std_logic                     := '0';             --                       reset.reset_n
		led_pio_external_connection_export : out   std_logic_vector(7 downto 0);                     -- led_pio_external_connection.export
		sdram_wire_addr                    : out   std_logic_vector(11 downto 0);                    --                  sdram_wire.addr
		sdram_wire_ba                      : out   std_logic_vector(1 downto 0);                     --                            .ba
		sdram_wire_cas_n                   : out   std_logic;                                        --                            .cas_n
		sdram_wire_cke                     : out   std_logic;                                        --                            .cke
		sdram_wire_cs_n                    : out   std_logic;                                        --                            .cs_n
		sdram_wire_dq                      : inout std_logic_vector(15 downto 0) := (others => '0'); --                            .dq
		sdram_wire_dqm                     : out   std_logic_vector(1 downto 0);                     --                            .dqm
		sdram_wire_ras_n                   : out   std_logic;                                        --                            .ras_n
		sdram_wire_we_n                    : out   std_logic                                         --                            .we_n
	);
end entity first_nios2_system;

architecture rtl of first_nios2_system is
	component first_nios2_system_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			M_ci_multi_done                       : in  std_logic                     := 'X';             -- done
			M_ci_multi_result                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_result
			M_ci_multi_a                          : out std_logic_vector(4 downto 0);                     -- multi_a
			M_ci_multi_b                          : out std_logic_vector(4 downto 0);                     -- multi_b
			M_ci_multi_c                          : out std_logic_vector(4 downto 0);                     -- multi_c
			M_ci_multi_clk_en                     : out std_logic;                                        -- clk_en
			A_ci_multi_clock                      : out std_logic;                                        -- clk
			A_ci_multi_reset                      : out std_logic;                                        -- reset
			A_ci_multi_reset_req                  : out std_logic;                                        -- reset_req
			M_ci_multi_dataa                      : out std_logic_vector(31 downto 0);                    -- multi_dataa
			M_ci_multi_datab                      : out std_logic_vector(31 downto 0);                    -- multi_datab
			M_ci_multi_n                          : out std_logic_vector(7 downto 0);                     -- multi_n
			M_ci_multi_readra                     : out std_logic;                                        -- multi_readra
			M_ci_multi_readrb                     : out std_logic;                                        -- multi_readrb
			M_ci_multi_start                      : out std_logic;                                        -- start
			M_ci_multi_writerc                    : out std_logic                                         -- multi_writerc
		);
	end component first_nios2_system_cpu;

	component first_nios2_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component first_nios2_system_jtag_uart;

	component first_nios2_system_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component first_nios2_system_sys_clk_timer;

	component first_nios2_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component first_nios2_system_sysid;

	component first_nios2_system_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component first_nios2_system_led_pio;

	component first_nios2_system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component first_nios2_system_sdram;

	component fp_mult is
		port (
			result : out std_logic_vector(31 downto 0);                    -- result
			clk    : in  std_logic                     := 'X';             -- clk
			start  : in  std_logic                     := 'X';             -- start
			done   : out std_logic;                                        -- done
			reset  : in  std_logic                     := 'X';             -- reset
			data   : in  std_logic_vector(31 downto 0) := (others => 'X')  -- dataa
		);
	end component fp_mult;

	component first_nios2_system_cpu_custom_instruction_master_translator is
		port (
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_c
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0)                      -- c
		);
	end component first_nios2_system_cpu_custom_instruction_master_translator;

	component first_nios2_system_cpu_custom_instruction_master_multi_xconnect is
		port (
			ci_slave_dataa       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result      : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra      : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb      : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc     : in  std_logic                     := 'X';             -- writerc
			ci_slave_a           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c           : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus     : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk         : in  std_logic                     := 'X';             -- clk
			ci_slave_reset       : in  std_logic                     := 'X';             -- reset
			ci_slave_clken       : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req   : in  std_logic                     := 'X';             -- reset_req
			ci_slave_start       : in  std_logic                     := 'X';             -- start
			ci_slave_done        : out std_logic;                                        -- done
			ci_master0_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra    : out std_logic;                                        -- readra
			ci_master0_readrb    : out std_logic;                                        -- readrb
			ci_master0_writerc   : out std_logic;                                        -- writerc
			ci_master0_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus   : out std_logic;                                        -- estatus
			ci_master0_clk       : out std_logic;                                        -- clk
			ci_master0_reset     : out std_logic;                                        -- reset
			ci_master0_clken     : out std_logic;                                        -- clk_en
			ci_master0_reset_req : out std_logic;                                        -- reset_req
			ci_master0_start     : out std_logic;                                        -- start
			ci_master0_done      : in  std_logic                     := 'X'              -- done
		);
	end component first_nios2_system_cpu_custom_instruction_master_multi_xconnect;

	component first_nios2_system_cpu_custom_instruction_master_multi_slave_translator0 is
		port (
			ci_slave_dataa     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result    : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra    : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb    : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc   : in  std_logic                     := 'X';             -- writerc
			ci_slave_a         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c         : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus   : in  std_logic                     := 'X';             -- estatus
			ci_slave_clk       : in  std_logic                     := 'X';             -- clk
			ci_slave_clken     : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req : in  std_logic                     := 'X';             -- reset_req
			ci_slave_reset     : in  std_logic                     := 'X';             -- reset
			ci_slave_start     : in  std_logic                     := 'X';             -- start
			ci_slave_done      : out std_logic;                                        -- done
			ci_master_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_clk      : out std_logic;                                        -- clk
			ci_master_clken    : out std_logic;                                        -- clk_en
			ci_master_reset    : out std_logic;                                        -- reset
			ci_master_start    : out std_logic;                                        -- start
			ci_master_done     : in  std_logic                     := 'X'              -- done
		);
	end component first_nios2_system_cpu_custom_instruction_master_multi_slave_translator0;

	component first_nios2_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                           : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                 : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address          : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			cpu_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write             : out std_logic;                                        -- write
			cpu_jtag_debug_module_read              : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			led_pio_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                        : out std_logic;                                        -- write
			led_pio_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                   : out std_logic;                                        -- chipselect
			sdram_s1_address                        : out std_logic_vector(21 downto 0);                    -- address
			sdram_s1_write                          : out std_logic;                                        -- write
			sdram_s1_read                           : out std_logic;                                        -- read
			sdram_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                     : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                  : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                     : out std_logic;                                        -- chipselect
			sys_clk_timer_s1_address                : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                  : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata              : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect             : out std_logic;                                        -- chipselect
			sysid_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component first_nios2_system_mm_interconnect_0;

	component first_nios2_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component first_nios2_system_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_custom_instruction_master_multi_readra                             : std_logic;                     -- cpu:M_ci_multi_readra -> cpu_custom_instruction_master_translator:ci_slave_multi_readra
	signal cpu_custom_instruction_master_multi_readrb                             : std_logic;                     -- cpu:M_ci_multi_readrb -> cpu_custom_instruction_master_translator:ci_slave_multi_readrb
	signal cpu_custom_instruction_master_multi_n                                  : std_logic_vector(7 downto 0);  -- cpu:M_ci_multi_n -> cpu_custom_instruction_master_translator:ci_slave_multi_n
	signal cpu_custom_instruction_master_done                                     : std_logic;                     -- cpu_custom_instruction_master_translator:ci_slave_multi_done -> cpu:M_ci_multi_done
	signal cpu_custom_instruction_master_clk_en                                   : std_logic;                     -- cpu:M_ci_multi_clk_en -> cpu_custom_instruction_master_translator:ci_slave_multi_clken
	signal cpu_custom_instruction_master_multi_writerc                            : std_logic;                     -- cpu:M_ci_multi_writerc -> cpu_custom_instruction_master_translator:ci_slave_multi_writerc
	signal cpu_custom_instruction_master_multi_result                             : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:ci_slave_multi_result -> cpu:M_ci_multi_result
	signal cpu_custom_instruction_master_clk                                      : std_logic;                     -- cpu:A_ci_multi_clock -> cpu_custom_instruction_master_translator:ci_slave_multi_clk
	signal cpu_custom_instruction_master_reset_req                                : std_logic;                     -- cpu:A_ci_multi_reset_req -> cpu_custom_instruction_master_translator:ci_slave_multi_reset_req
	signal cpu_custom_instruction_master_multi_c                                  : std_logic_vector(4 downto 0);  -- cpu:M_ci_multi_c -> cpu_custom_instruction_master_translator:ci_slave_multi_c
	signal cpu_custom_instruction_master_multi_b                                  : std_logic_vector(4 downto 0);  -- cpu:M_ci_multi_b -> cpu_custom_instruction_master_translator:ci_slave_multi_b
	signal cpu_custom_instruction_master_multi_a                                  : std_logic_vector(4 downto 0);  -- cpu:M_ci_multi_a -> cpu_custom_instruction_master_translator:ci_slave_multi_a
	signal cpu_custom_instruction_master_multi_dataa                              : std_logic_vector(31 downto 0); -- cpu:M_ci_multi_dataa -> cpu_custom_instruction_master_translator:ci_slave_multi_dataa
	signal cpu_custom_instruction_master_start                                    : std_logic;                     -- cpu:M_ci_multi_start -> cpu_custom_instruction_master_translator:ci_slave_multi_start
	signal cpu_custom_instruction_master_multi_datab                              : std_logic_vector(31 downto 0); -- cpu:M_ci_multi_datab -> cpu_custom_instruction_master_translator:ci_slave_multi_datab
	signal cpu_custom_instruction_master_reset                                    : std_logic;                     -- cpu:A_ci_multi_reset -> cpu_custom_instruction_master_translator:ci_slave_multi_reset
	signal cpu_custom_instruction_master_translator_multi_ci_master_result        : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:multi_ci_master_result
	signal cpu_custom_instruction_master_translator_multi_ci_master_b             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_b -> cpu_custom_instruction_master_multi_xconnect:ci_slave_b
	signal cpu_custom_instruction_master_translator_multi_ci_master_c             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_c -> cpu_custom_instruction_master_multi_xconnect:ci_slave_c
	signal cpu_custom_instruction_master_translator_multi_ci_master_a             : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_a -> cpu_custom_instruction_master_multi_xconnect:ci_slave_a
	signal cpu_custom_instruction_master_translator_multi_ci_master_clk_en        : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_clken -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clken
	signal cpu_custom_instruction_master_translator_multi_ci_master_done          : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_custom_instruction_master_translator:multi_ci_master_done
	signal cpu_custom_instruction_master_translator_multi_ci_master_n             : std_logic_vector(7 downto 0);  -- cpu_custom_instruction_master_translator:multi_ci_master_n -> cpu_custom_instruction_master_multi_xconnect:ci_slave_n
	signal cpu_custom_instruction_master_translator_multi_ci_master_writerc       : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_custom_instruction_master_multi_xconnect:ci_slave_writerc
	signal cpu_custom_instruction_master_translator_multi_ci_master_clk           : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_clk -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clk
	signal cpu_custom_instruction_master_translator_multi_ci_master_reset_req     : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	signal cpu_custom_instruction_master_translator_multi_ci_master_start         : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_start -> cpu_custom_instruction_master_multi_xconnect:ci_slave_start
	signal cpu_custom_instruction_master_translator_multi_ci_master_dataa         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_custom_instruction_master_multi_xconnect:ci_slave_dataa
	signal cpu_custom_instruction_master_translator_multi_ci_master_readra        : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_readra -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readra
	signal cpu_custom_instruction_master_translator_multi_ci_master_reset         : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_reset -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset
	signal cpu_custom_instruction_master_translator_multi_ci_master_datab         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_translator:multi_ci_master_datab -> cpu_custom_instruction_master_multi_xconnect:ci_slave_datab
	signal cpu_custom_instruction_master_translator_multi_ci_master_readrb        : std_logic;                     -- cpu_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readrb
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_multi_xconnect:ci_master0_result
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_b
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_c
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_done           : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_custom_instruction_master_multi_xconnect:ci_master0_done
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en         : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_a
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- cpu_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_n
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc        : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_clk            : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req      : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_start          : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_start
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_readra         : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_reset          : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb         : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	signal cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus        : std_logic;                     -- cpu_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- fp_mult_0:result -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_result
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_start  : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_start -> fp_mult_0:start
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> fp_mult_0:data
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_done   : std_logic;                     -- fp_mult_0:done -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_done
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset  : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset -> fp_mult_0:reset
	signal cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk    : std_logic;                     -- cpu_custom_instruction_master_multi_slave_translator0:ci_master_clk -> fp_mult_0:clk
	signal cpu_instruction_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                         : std_logic_vector(24 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                            : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_0_led_pio_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_0_led_pio_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_write                                     : std_logic;                     -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_readdata                                  : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_sys_clk_timer_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_write                               : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                            : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                 : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_writedata                                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_sdram_s1_address                                     : std_logic_vector(21 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_write                                       : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_read                                        : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_readdata                                    : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_readdatavalid                               : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_byteenable                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sysid_control_slave_address                          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_sysid_control_slave_readdata                         : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest                    : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal mm_interconnect_0_cpu_jtag_debug_module_address                        : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_write                          : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_read                           : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata                       : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess                    : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal cpu_data_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                              : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_data_master_address                                                : std_logic_vector(24 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_write                                                  : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_read                                                   : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_debugaccess                                            : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_byteenable                                             : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest              : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect               : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                    : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                     : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                 : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal irq_mapper_receiver0_irq                                               : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                               : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal rst_controller_reset_out_reset                                         : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                     : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                                : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                              : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv           : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal rst_controller_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n, led_pio:reset_n, sdram:reset_n, sys_clk_timer:reset_n, sysid:reset_n]

begin

	cpu : component first_nios2_system_cpu
		port map (
			clk                                   => clk_clk,                                             --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,   --                          .writedata
			M_ci_multi_done                       => cpu_custom_instruction_master_done,                  -- custom_instruction_master.done
			M_ci_multi_result                     => cpu_custom_instruction_master_multi_result,          --                          .multi_result
			M_ci_multi_a                          => cpu_custom_instruction_master_multi_a,               --                          .multi_a
			M_ci_multi_b                          => cpu_custom_instruction_master_multi_b,               --                          .multi_b
			M_ci_multi_c                          => cpu_custom_instruction_master_multi_c,               --                          .multi_c
			M_ci_multi_clk_en                     => cpu_custom_instruction_master_clk_en,                --                          .clk_en
			A_ci_multi_clock                      => cpu_custom_instruction_master_clk,                   --                          .clk
			A_ci_multi_reset                      => cpu_custom_instruction_master_reset,                 --                          .reset
			A_ci_multi_reset_req                  => cpu_custom_instruction_master_reset_req,             --                          .reset_req
			M_ci_multi_dataa                      => cpu_custom_instruction_master_multi_dataa,           --                          .multi_dataa
			M_ci_multi_datab                      => cpu_custom_instruction_master_multi_datab,           --                          .multi_datab
			M_ci_multi_n                          => cpu_custom_instruction_master_multi_n,               --                          .multi_n
			M_ci_multi_readra                     => cpu_custom_instruction_master_multi_readra,          --                          .multi_readra
			M_ci_multi_readrb                     => cpu_custom_instruction_master_multi_readrb,          --                          .multi_readrb
			M_ci_multi_start                      => cpu_custom_instruction_master_start,                 --                          .start
			M_ci_multi_writerc                    => cpu_custom_instruction_master_multi_writerc          --                          .multi_writerc
		);

	jtag_uart : component first_nios2_system_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	sys_clk_timer : component first_nios2_system_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                            --   irq.irq
		);

	sysid : component first_nios2_system_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	led_pio : component first_nios2_system_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	sdram : component first_nios2_system_sdram
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	fp_mult_0 : component fp_mult
		port map (
			result => cpu_custom_instruction_master_multi_slave_translator0_ci_master_result, -- fp_mult.result
			clk    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --        .clk
			start  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_start,  --        .start
			done   => cpu_custom_instruction_master_multi_slave_translator0_ci_master_done,   --        .done
			reset  => cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --        .reset
			data   => cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa   --        .dataa
		);

	cpu_custom_instruction_master_translator : component first_nios2_system_cpu_custom_instruction_master_translator
		port map (
			ci_slave_result           => open,                                                               --        ci_slave.result
			ci_slave_multi_clk        => cpu_custom_instruction_master_clk,                                  --                .clk
			ci_slave_multi_reset      => cpu_custom_instruction_master_reset,                                --                .reset
			ci_slave_multi_clken      => cpu_custom_instruction_master_clk_en,                               --                .clk_en
			ci_slave_multi_reset_req  => cpu_custom_instruction_master_reset_req,                            --                .reset_req
			ci_slave_multi_start      => cpu_custom_instruction_master_start,                                --                .start
			ci_slave_multi_done       => cpu_custom_instruction_master_done,                                 --                .done
			ci_slave_multi_dataa      => cpu_custom_instruction_master_multi_dataa,                          --                .multi_dataa
			ci_slave_multi_datab      => cpu_custom_instruction_master_multi_datab,                          --                .multi_datab
			ci_slave_multi_result     => cpu_custom_instruction_master_multi_result,                         --                .multi_result
			ci_slave_multi_n          => cpu_custom_instruction_master_multi_n,                              --                .multi_n
			ci_slave_multi_readra     => cpu_custom_instruction_master_multi_readra,                         --                .multi_readra
			ci_slave_multi_readrb     => cpu_custom_instruction_master_multi_readrb,                         --                .multi_readrb
			ci_slave_multi_writerc    => cpu_custom_instruction_master_multi_writerc,                        --                .multi_writerc
			ci_slave_multi_a          => cpu_custom_instruction_master_multi_a,                              --                .multi_a
			ci_slave_multi_b          => cpu_custom_instruction_master_multi_b,                              --                .multi_b
			ci_slave_multi_c          => cpu_custom_instruction_master_multi_c,                              --                .multi_c
			comb_ci_master_result     => open,                                                               --  comb_ci_master.result
			multi_ci_master_clk       => cpu_custom_instruction_master_translator_multi_ci_master_clk,       -- multi_ci_master.clk
			multi_ci_master_reset     => cpu_custom_instruction_master_translator_multi_ci_master_reset,     --                .reset
			multi_ci_master_clken     => cpu_custom_instruction_master_translator_multi_ci_master_clk_en,    --                .clk_en
			multi_ci_master_reset_req => cpu_custom_instruction_master_translator_multi_ci_master_reset_req, --                .reset_req
			multi_ci_master_start     => cpu_custom_instruction_master_translator_multi_ci_master_start,     --                .start
			multi_ci_master_done      => cpu_custom_instruction_master_translator_multi_ci_master_done,      --                .done
			multi_ci_master_dataa     => cpu_custom_instruction_master_translator_multi_ci_master_dataa,     --                .dataa
			multi_ci_master_datab     => cpu_custom_instruction_master_translator_multi_ci_master_datab,     --                .datab
			multi_ci_master_result    => cpu_custom_instruction_master_translator_multi_ci_master_result,    --                .result
			multi_ci_master_n         => cpu_custom_instruction_master_translator_multi_ci_master_n,         --                .n
			multi_ci_master_readra    => cpu_custom_instruction_master_translator_multi_ci_master_readra,    --                .readra
			multi_ci_master_readrb    => cpu_custom_instruction_master_translator_multi_ci_master_readrb,    --                .readrb
			multi_ci_master_writerc   => cpu_custom_instruction_master_translator_multi_ci_master_writerc,   --                .writerc
			multi_ci_master_a         => cpu_custom_instruction_master_translator_multi_ci_master_a,         --                .a
			multi_ci_master_b         => cpu_custom_instruction_master_translator_multi_ci_master_b,         --                .b
			multi_ci_master_c         => cpu_custom_instruction_master_translator_multi_ci_master_c          --                .c
		);

	cpu_custom_instruction_master_multi_xconnect : component first_nios2_system_cpu_custom_instruction_master_multi_xconnect
		port map (
			ci_slave_dataa       => cpu_custom_instruction_master_translator_multi_ci_master_dataa,     --   ci_slave.dataa
			ci_slave_datab       => cpu_custom_instruction_master_translator_multi_ci_master_datab,     --           .datab
			ci_slave_result      => cpu_custom_instruction_master_translator_multi_ci_master_result,    --           .result
			ci_slave_n           => cpu_custom_instruction_master_translator_multi_ci_master_n,         --           .n
			ci_slave_readra      => cpu_custom_instruction_master_translator_multi_ci_master_readra,    --           .readra
			ci_slave_readrb      => cpu_custom_instruction_master_translator_multi_ci_master_readrb,    --           .readrb
			ci_slave_writerc     => cpu_custom_instruction_master_translator_multi_ci_master_writerc,   --           .writerc
			ci_slave_a           => cpu_custom_instruction_master_translator_multi_ci_master_a,         --           .a
			ci_slave_b           => cpu_custom_instruction_master_translator_multi_ci_master_b,         --           .b
			ci_slave_c           => cpu_custom_instruction_master_translator_multi_ci_master_c,         --           .c
			ci_slave_ipending    => open,                                                               --           .ipending
			ci_slave_estatus     => open,                                                               --           .estatus
			ci_slave_clk         => cpu_custom_instruction_master_translator_multi_ci_master_clk,       --           .clk
			ci_slave_reset       => cpu_custom_instruction_master_translator_multi_ci_master_reset,     --           .reset
			ci_slave_clken       => cpu_custom_instruction_master_translator_multi_ci_master_clk_en,    --           .clk_en
			ci_slave_reset_req   => cpu_custom_instruction_master_translator_multi_ci_master_reset_req, --           .reset_req
			ci_slave_start       => cpu_custom_instruction_master_translator_multi_ci_master_start,     --           .start
			ci_slave_done        => cpu_custom_instruction_master_translator_multi_ci_master_done,      --           .done
			ci_master0_dataa     => cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa,      -- ci_master0.dataa
			ci_master0_datab     => cpu_custom_instruction_master_multi_xconnect_ci_master0_datab,      --           .datab
			ci_master0_result    => cpu_custom_instruction_master_multi_xconnect_ci_master0_result,     --           .result
			ci_master0_n         => cpu_custom_instruction_master_multi_xconnect_ci_master0_n,          --           .n
			ci_master0_readra    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readra,     --           .readra
			ci_master0_readrb    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb,     --           .readrb
			ci_master0_writerc   => cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc,    --           .writerc
			ci_master0_a         => cpu_custom_instruction_master_multi_xconnect_ci_master0_a,          --           .a
			ci_master0_b         => cpu_custom_instruction_master_multi_xconnect_ci_master0_b,          --           .b
			ci_master0_c         => cpu_custom_instruction_master_multi_xconnect_ci_master0_c,          --           .c
			ci_master0_ipending  => cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending,   --           .ipending
			ci_master0_estatus   => cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus,    --           .estatus
			ci_master0_clk       => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk,        --           .clk
			ci_master0_reset     => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset,      --           .reset
			ci_master0_clken     => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en,     --           .clk_en
			ci_master0_reset_req => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req,  --           .reset_req
			ci_master0_start     => cpu_custom_instruction_master_multi_xconnect_ci_master0_start,      --           .start
			ci_master0_done      => cpu_custom_instruction_master_multi_xconnect_ci_master0_done        --           .done
		);

	cpu_custom_instruction_master_multi_slave_translator0 : component first_nios2_system_cpu_custom_instruction_master_multi_slave_translator0
		port map (
			ci_slave_dataa     => cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab     => cpu_custom_instruction_master_multi_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result    => cpu_custom_instruction_master_multi_xconnect_ci_master0_result,         --          .result
			ci_slave_n         => cpu_custom_instruction_master_multi_xconnect_ci_master0_n,              --          .n
			ci_slave_readra    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb    => cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc   => cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a         => cpu_custom_instruction_master_multi_xconnect_ci_master0_a,              --          .a
			ci_slave_b         => cpu_custom_instruction_master_multi_xconnect_ci_master0_b,              --          .b
			ci_slave_c         => cpu_custom_instruction_master_multi_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending  => cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus   => cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus,        --          .estatus
			ci_slave_clk       => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk,            --          .clk
			ci_slave_clken     => cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en,         --          .clk_en
			ci_slave_reset_req => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req,      --          .reset_req
			ci_slave_reset     => cpu_custom_instruction_master_multi_xconnect_ci_master0_reset,          --          .reset
			ci_slave_start     => cpu_custom_instruction_master_multi_xconnect_ci_master0_start,          --          .start
			ci_slave_done      => cpu_custom_instruction_master_multi_xconnect_ci_master0_done,           --          .done
			ci_master_dataa    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_result   => cpu_custom_instruction_master_multi_slave_translator0_ci_master_result, --          .result
			ci_master_clk      => cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk,    --          .clk
			ci_master_clken    => open,                                                                   --          .clk_en
			ci_master_reset    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset,  --          .reset
			ci_master_start    => cpu_custom_instruction_master_multi_slave_translator0_ci_master_start,  --          .start
			ci_master_done     => cpu_custom_instruction_master_multi_slave_translator0_ci_master_done    --          .done
		);

	mm_interconnect_0 : component first_nios2_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                           => clk_clk,                                                   --                         clk_0_clk.clk
			cpu_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- cpu_reset_n_reset_bridge_in_reset.reset
			cpu_data_master_address                 => cpu_data_master_address,                                   --                   cpu_data_master.address
			cpu_data_master_waitrequest             => cpu_data_master_waitrequest,                               --                                  .waitrequest
			cpu_data_master_byteenable              => cpu_data_master_byteenable,                                --                                  .byteenable
			cpu_data_master_read                    => cpu_data_master_read,                                      --                                  .read
			cpu_data_master_readdata                => cpu_data_master_readdata,                                  --                                  .readdata
			cpu_data_master_write                   => cpu_data_master_write,                                     --                                  .write
			cpu_data_master_writedata               => cpu_data_master_writedata,                                 --                                  .writedata
			cpu_data_master_debugaccess             => cpu_data_master_debugaccess,                               --                                  .debugaccess
			cpu_instruction_master_address          => cpu_instruction_master_address,                            --            cpu_instruction_master.address
			cpu_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                        --                                  .waitrequest
			cpu_instruction_master_read             => cpu_instruction_master_read,                               --                                  .read
			cpu_instruction_master_readdata         => cpu_instruction_master_readdata,                           --                                  .readdata
			cpu_instruction_master_readdatavalid    => cpu_instruction_master_readdatavalid,                      --                                  .readdatavalid
			cpu_jtag_debug_module_address           => mm_interconnect_0_cpu_jtag_debug_module_address,           --             cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write             => mm_interconnect_0_cpu_jtag_debug_module_write,             --                                  .write
			cpu_jtag_debug_module_read              => mm_interconnect_0_cpu_jtag_debug_module_read,              --                                  .read
			cpu_jtag_debug_module_readdata          => mm_interconnect_0_cpu_jtag_debug_module_readdata,          --                                  .readdata
			cpu_jtag_debug_module_writedata         => mm_interconnect_0_cpu_jtag_debug_module_writedata,         --                                  .writedata
			cpu_jtag_debug_module_byteenable        => mm_interconnect_0_cpu_jtag_debug_module_byteenable,        --                                  .byteenable
			cpu_jtag_debug_module_waitrequest       => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,       --                                  .waitrequest
			cpu_jtag_debug_module_debugaccess       => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,       --                                  .debugaccess
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --       jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                  .chipselect
			led_pio_s1_address                      => mm_interconnect_0_led_pio_s1_address,                      --                        led_pio_s1.address
			led_pio_s1_write                        => mm_interconnect_0_led_pio_s1_write,                        --                                  .write
			led_pio_s1_readdata                     => mm_interconnect_0_led_pio_s1_readdata,                     --                                  .readdata
			led_pio_s1_writedata                    => mm_interconnect_0_led_pio_s1_writedata,                    --                                  .writedata
			led_pio_s1_chipselect                   => mm_interconnect_0_led_pio_s1_chipselect,                   --                                  .chipselect
			sdram_s1_address                        => mm_interconnect_0_sdram_s1_address,                        --                          sdram_s1.address
			sdram_s1_write                          => mm_interconnect_0_sdram_s1_write,                          --                                  .write
			sdram_s1_read                           => mm_interconnect_0_sdram_s1_read,                           --                                  .read
			sdram_s1_readdata                       => mm_interconnect_0_sdram_s1_readdata,                       --                                  .readdata
			sdram_s1_writedata                      => mm_interconnect_0_sdram_s1_writedata,                      --                                  .writedata
			sdram_s1_byteenable                     => mm_interconnect_0_sdram_s1_byteenable,                     --                                  .byteenable
			sdram_s1_readdatavalid                  => mm_interconnect_0_sdram_s1_readdatavalid,                  --                                  .readdatavalid
			sdram_s1_waitrequest                    => mm_interconnect_0_sdram_s1_waitrequest,                    --                                  .waitrequest
			sdram_s1_chipselect                     => mm_interconnect_0_sdram_s1_chipselect,                     --                                  .chipselect
			sys_clk_timer_s1_address                => mm_interconnect_0_sys_clk_timer_s1_address,                --                  sys_clk_timer_s1.address
			sys_clk_timer_s1_write                  => mm_interconnect_0_sys_clk_timer_s1_write,                  --                                  .write
			sys_clk_timer_s1_readdata               => mm_interconnect_0_sys_clk_timer_s1_readdata,               --                                  .readdata
			sys_clk_timer_s1_writedata              => mm_interconnect_0_sys_clk_timer_s1_writedata,              --                                  .writedata
			sys_clk_timer_s1_chipselect             => mm_interconnect_0_sys_clk_timer_s1_chipselect,             --                                  .chipselect
			sysid_control_slave_address             => mm_interconnect_0_sysid_control_slave_address,             --               sysid_control_slave.address
			sysid_control_slave_readdata            => mm_interconnect_0_sysid_control_slave_readdata             --                                  .readdata
		);

	irq_mapper : component first_nios2_system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of first_nios2_system
