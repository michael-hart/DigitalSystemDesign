// first_nios2_system.v

// Generated using ACDS version 13.1 162 at 2016.03.04.13:55:27

`timescale 1 ps / 1 ps
module first_nios2_system (
		input  wire        clk_clk,                            //                         clk.clk
		input  wire        reset_reset_n,                      //                       reset.reset_n
		output wire [7:0]  led_pio_external_connection_export, // led_pio_external_connection.export
		output wire [11:0] sdram_wire_addr,                    //                  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                      //                            .ba
		output wire        sdram_wire_cas_n,                   //                            .cas_n
		output wire        sdram_wire_cke,                     //                            .cke
		output wire        sdram_wire_cs_n,                    //                            .cs_n
		inout  wire [15:0] sdram_wire_dq,                      //                            .dq
		output wire [1:0]  sdram_wire_dqm,                     //                            .dqm
		output wire        sdram_wire_ras_n,                   //                            .ras_n
		output wire        sdram_wire_we_n                     //                            .we_n
	);

	wire         cpu_custom_instruction_master_multi_readra;                             // cpu:M_ci_multi_readra -> cpu_custom_instruction_master_translator:ci_slave_multi_readra
	wire         cpu_custom_instruction_master_multi_readrb;                             // cpu:M_ci_multi_readrb -> cpu_custom_instruction_master_translator:ci_slave_multi_readrb
	wire   [7:0] cpu_custom_instruction_master_multi_n;                                  // cpu:M_ci_multi_n -> cpu_custom_instruction_master_translator:ci_slave_multi_n
	wire         cpu_custom_instruction_master_done;                                     // cpu_custom_instruction_master_translator:ci_slave_multi_done -> cpu:M_ci_multi_done
	wire         cpu_custom_instruction_master_clk_en;                                   // cpu:M_ci_multi_clk_en -> cpu_custom_instruction_master_translator:ci_slave_multi_clken
	wire         cpu_custom_instruction_master_multi_writerc;                            // cpu:M_ci_multi_writerc -> cpu_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] cpu_custom_instruction_master_multi_result;                             // cpu_custom_instruction_master_translator:ci_slave_multi_result -> cpu:M_ci_multi_result
	wire         cpu_custom_instruction_master_clk;                                      // cpu:A_ci_multi_clock -> cpu_custom_instruction_master_translator:ci_slave_multi_clk
	wire         cpu_custom_instruction_master_reset_req;                                // cpu:A_ci_multi_reset_req -> cpu_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] cpu_custom_instruction_master_multi_c;                                  // cpu:M_ci_multi_c -> cpu_custom_instruction_master_translator:ci_slave_multi_c
	wire   [4:0] cpu_custom_instruction_master_multi_b;                                  // cpu:M_ci_multi_b -> cpu_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] cpu_custom_instruction_master_multi_a;                                  // cpu:M_ci_multi_a -> cpu_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] cpu_custom_instruction_master_multi_dataa;                              // cpu:M_ci_multi_dataa -> cpu_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         cpu_custom_instruction_master_start;                                    // cpu:M_ci_multi_start -> cpu_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] cpu_custom_instruction_master_multi_datab;                              // cpu:M_ci_multi_datab -> cpu_custom_instruction_master_translator:ci_slave_multi_datab
	wire         cpu_custom_instruction_master_reset;                                    // cpu:A_ci_multi_reset -> cpu_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_result;        // cpu_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_b;             // cpu_custom_instruction_master_translator:multi_ci_master_b -> cpu_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_c;             // cpu_custom_instruction_master_translator:multi_ci_master_c -> cpu_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_a;             // cpu_custom_instruction_master_translator:multi_ci_master_a -> cpu_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         cpu_custom_instruction_master_translator_multi_ci_master_clk_en;        // cpu_custom_instruction_master_translator:multi_ci_master_clken -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         cpu_custom_instruction_master_translator_multi_ci_master_done;          // cpu_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu_custom_instruction_master_translator_multi_ci_master_n;             // cpu_custom_instruction_master_translator:multi_ci_master_n -> cpu_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         cpu_custom_instruction_master_translator_multi_ci_master_writerc;       // cpu_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu_custom_instruction_master_translator_multi_ci_master_clk;           // cpu_custom_instruction_master_translator:multi_ci_master_clk -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu_custom_instruction_master_translator_multi_ci_master_reset_req;     // cpu_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu_custom_instruction_master_translator_multi_ci_master_start;         // cpu_custom_instruction_master_translator:multi_ci_master_start -> cpu_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_dataa;         // cpu_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu_custom_instruction_master_translator_multi_ci_master_readra;        // cpu_custom_instruction_master_translator:multi_ci_master_readra -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         cpu_custom_instruction_master_translator_multi_ci_master_reset;         // cpu_custom_instruction_master_translator:multi_ci_master_reset -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_datab;         // cpu_custom_instruction_master_translator:multi_ci_master_datab -> cpu_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         cpu_custom_instruction_master_translator_multi_ci_master_readrb;        // cpu_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_result;         // cpu_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_b;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_c;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_done;           // cpu_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // cpu_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_a;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_n;              // cpu_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // cpu_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // cpu_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_clk;            // cpu_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // cpu_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_start;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_readra;         // cpu_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_reset;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_datab;          // cpu_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // cpu_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // cpu_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_result; // fp_mult_0:result -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_start;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_start -> fp_mult_0:start
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> fp_mult_0:dataa
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_done;   // fp_mult_0:done -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_n;      // cpu_custom_instruction_master_multi_slave_translator0:ci_master_n -> fp_mult_0:opcode
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset -> fp_mult_0:resetn
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // cpu_custom_instruction_master_multi_slave_translator0:ci_master_datab -> fp_mult_0:datab
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // cpu_custom_instruction_master_multi_slave_translator0:ci_master_clk -> fp_mult_0:clk
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                          // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                         // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;              // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                 // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                           // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                             // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;                          // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                               // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                            // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                                 // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                                   // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_chipselect;                                // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire         mm_interconnect_0_led_pio_s1_write;                                     // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                                  // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                    // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                      // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                        // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                          // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                           // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                       // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                    // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                     // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         cpu_data_master_waitrequest;                                            // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                              // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [24:0] cpu_data_master_address;                                                // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                                  // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                                   // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                               // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                            // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                             // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_instruction_master_waitrequest;                                     // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [24:0] cpu_instruction_master_address;                                         // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                            // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                        // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                                   // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                 // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                   // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                                     // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                  // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                       // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                        // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                    // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                               // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                  // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         irq_mapper_receiver0_irq;                                               // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                               // sys_clk_timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                                          // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, led_pio:reset_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]

	first_nios2_system_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                    //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.M_ci_multi_done                       (cpu_custom_instruction_master_done),                  // custom_instruction_master.done
		.M_ci_multi_result                     (cpu_custom_instruction_master_multi_result),          //                          .multi_result
		.M_ci_multi_a                          (cpu_custom_instruction_master_multi_a),               //                          .multi_a
		.M_ci_multi_b                          (cpu_custom_instruction_master_multi_b),               //                          .multi_b
		.M_ci_multi_c                          (cpu_custom_instruction_master_multi_c),               //                          .multi_c
		.M_ci_multi_clk_en                     (cpu_custom_instruction_master_clk_en),                //                          .clk_en
		.A_ci_multi_clock                      (cpu_custom_instruction_master_clk),                   //                          .clk
		.A_ci_multi_reset                      (cpu_custom_instruction_master_reset),                 //                          .reset
		.A_ci_multi_reset_req                  (cpu_custom_instruction_master_reset_req),             //                          .reset_req
		.M_ci_multi_dataa                      (cpu_custom_instruction_master_multi_dataa),           //                          .multi_dataa
		.M_ci_multi_datab                      (cpu_custom_instruction_master_multi_datab),           //                          .multi_datab
		.M_ci_multi_n                          (cpu_custom_instruction_master_multi_n),               //                          .multi_n
		.M_ci_multi_readra                     (cpu_custom_instruction_master_multi_readra),          //                          .multi_readra
		.M_ci_multi_readrb                     (cpu_custom_instruction_master_multi_readrb),          //                          .multi_readrb
		.M_ci_multi_start                      (cpu_custom_instruction_master_start),                 //                          .start
		.M_ci_multi_writerc                    (cpu_custom_instruction_master_multi_writerc)          //                          .multi_writerc
	);

	first_nios2_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	first_nios2_system_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                       //   irq.irq
	);

	first_nios2_system_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	first_nios2_system_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)       // external_connection.export
	);

	first_nios2_system_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	fp_mult fp_mult_0 (
		.opcode (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),      // fp_mult.n
		.dataa  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //        .dataa
		.datab  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //        .datab
		.result (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result), //        .result
		.clk    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //        .clk
		.start  (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),  //        .start
		.resetn (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //        .reset
		.done   (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done)    //        .done
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                   //        ci_slave.result
		.ci_slave_multi_clk        (cpu_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (cpu_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (cpu_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (cpu_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (cpu_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (cpu_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (cpu_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (cpu_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (cpu_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (cpu_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (cpu_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                   //  comb_ci_master.result
		.multi_ci_master_clk       (cpu_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_n                (8'b00000000),                                                        //     (terminated)
		.ci_slave_readra           (1'b0),                                                               //     (terminated)
		.ci_slave_readrb           (1'b0),                                                               //     (terminated)
		.ci_slave_writerc          (1'b0),                                                               //     (terminated)
		.ci_slave_a                (5'b00000),                                                           //     (terminated)
		.ci_slave_b                (5'b00000),                                                           //     (terminated)
		.ci_slave_c                (5'b00000),                                                           //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_estatus          (1'b0),                                                               //     (terminated)
		.comb_ci_master_dataa      (),                                                                   //     (terminated)
		.comb_ci_master_datab      (),                                                                   //     (terminated)
		.comb_ci_master_n          (),                                                                   //     (terminated)
		.comb_ci_master_readra     (),                                                                   //     (terminated)
		.comb_ci_master_readrb     (),                                                                   //     (terminated)
		.comb_ci_master_writerc    (),                                                                   //     (terminated)
		.comb_ci_master_a          (),                                                                   //     (terminated)
		.comb_ci_master_b          (),                                                                   //     (terminated)
		.comb_ci_master_c          (),                                                                   //     (terminated)
		.comb_ci_master_ipending   (),                                                                   //     (terminated)
		.comb_ci_master_estatus    ()                                                                    //     (terminated)
	);

	first_nios2_system_cpu_custom_instruction_master_multi_xconnect cpu_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                   //           .ipending
		.ci_slave_estatus     (),                                                                   //           .estatus
		.ci_slave_clk         (cpu_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (cpu_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (),                                                                       //          .clk_en
		.ci_master_reset     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                       // (terminated)
		.ci_master_readrb    (),                                                                       // (terminated)
		.ci_master_writerc   (),                                                                       // (terminated)
		.ci_master_a         (),                                                                       // (terminated)
		.ci_master_b         (),                                                                       // (terminated)
		.ci_master_c         (),                                                                       // (terminated)
		.ci_master_ipending  (),                                                                       // (terminated)
		.ci_master_estatus   (),                                                                       // (terminated)
		.ci_master_reset_req ()                                                                        // (terminated)
	);

	first_nios2_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                         clk_0_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                  .readdatavalid
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.led_pio_s1_address                      (mm_interconnect_0_led_pio_s1_address),                      //                        led_pio_s1.address
		.led_pio_s1_write                        (mm_interconnect_0_led_pio_s1_write),                        //                                  .write
		.led_pio_s1_readdata                     (mm_interconnect_0_led_pio_s1_readdata),                     //                                  .readdata
		.led_pio_s1_writedata                    (mm_interconnect_0_led_pio_s1_writedata),                    //                                  .writedata
		.led_pio_s1_chipselect                   (mm_interconnect_0_led_pio_s1_chipselect),                   //                                  .chipselect
		.sdram_s1_address                        (mm_interconnect_0_sdram_s1_address),                        //                          sdram_s1.address
		.sdram_s1_write                          (mm_interconnect_0_sdram_s1_write),                          //                                  .write
		.sdram_s1_read                           (mm_interconnect_0_sdram_s1_read),                           //                                  .read
		.sdram_s1_readdata                       (mm_interconnect_0_sdram_s1_readdata),                       //                                  .readdata
		.sdram_s1_writedata                      (mm_interconnect_0_sdram_s1_writedata),                      //                                  .writedata
		.sdram_s1_byteenable                     (mm_interconnect_0_sdram_s1_byteenable),                     //                                  .byteenable
		.sdram_s1_readdatavalid                  (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                  .readdatavalid
		.sdram_s1_waitrequest                    (mm_interconnect_0_sdram_s1_waitrequest),                    //                                  .waitrequest
		.sdram_s1_chipselect                     (mm_interconnect_0_sdram_s1_chipselect),                     //                                  .chipselect
		.sys_clk_timer_s1_address                (mm_interconnect_0_sys_clk_timer_s1_address),                //                  sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                  (mm_interconnect_0_sys_clk_timer_s1_write),                  //                                  .write
		.sys_clk_timer_s1_readdata               (mm_interconnect_0_sys_clk_timer_s1_readdata),               //                                  .readdata
		.sys_clk_timer_s1_writedata              (mm_interconnect_0_sys_clk_timer_s1_writedata),              //                                  .writedata
		.sys_clk_timer_s1_chipselect             (mm_interconnect_0_sys_clk_timer_s1_chipselect),             //                                  .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //               sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata)             //                                  .readdata
	);

	first_nios2_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
